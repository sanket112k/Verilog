module n_bit_bcd_adder_tb;
parameter N=2;
parameter B=N*$clog2(10);
reg [N*4-1:0]bcd_in1,bcd_in2;
reg cin;
wire cout;
wire [N*4-1:0]sum;
integer i1,j1,k1,i2,j2,k2;
reg [B+N*4:0]shift_reg1,shift_reg2;
n_bit_bcd_adder #(.N(N)) dut(bcd_in1,bcd_in2,cin,cout,sum);
initial begin
    cin=0;
    shift_reg1=0;
    for(k1=0;k1<=(2**B)-1;k1=k1+1) begin
        if(shift_reg1[B+N*4-1:B]!={N{4'h9}}) begin
            shift_reg1[B+N*4:B]=0;
            shift_reg1[B-1:0]=k1;
            for(i1=0;i1<B;i1=i1+1) begin
                for(j1=0;j1<B;j1=j1+1) begin
                    if(shift_reg1[B+j1*4 +: 4]>=5)
                        shift_reg1[B+j1*4 +: 4] = shift_reg1[B+j1*4 +: 4] + 3;
                end
                shift_reg1=shift_reg1<<1;
            end
            bcd_in1=shift_reg1[B+N*4-1:B];
            shift_reg2=0;
            for(k2=0;k2<=(2**B)-1;k2=k2+1) begin
                if(shift_reg2[B+N*4-1:B]!={N{4'h9}}) begin
                    shift_reg2[B+N*4:B]=0;
                    shift_reg2[B-1:0]=k2;
                    for(i2=0;i2<B;i2=i2+1) begin
                        for(j2=0;j2<B;j2=j2+1) begin
                            if(shift_reg2[B+j2*4 +: 4]>=5)
                                shift_reg2[B+j2*4 +: 4] = shift_reg2[B+j2*4 +: 4] + 3;
                        end
                        shift_reg2=shift_reg2<<1;
                    end
                    bcd_in2=shift_reg2[B+N*4-1:B];
                    #10;
                end
            end
            #10;
        end
    end
    $finish;
end
initial begin
    $monitor("bcd_in1=%b bcd_in2=%b cout=%b sum=%b",bcd_in1,bcd_in2,cout,sum);
end
endmodule


/*
* OUTPUT
* bcd_in1=00000000 bcd_in2=00000000 cout=0 sum=00000000
* bcd_in1=00000000 bcd_in2=00000001 cout=0 sum=00000001
* bcd_in1=00000000 bcd_in2=00000010 cout=0 sum=00000010
* bcd_in1=00000000 bcd_in2=00000011 cout=0 sum=00000011
* bcd_in1=00000000 bcd_in2=00000100 cout=0 sum=00000100
* bcd_in1=00000000 bcd_in2=00000101 cout=0 sum=00000101
* bcd_in1=00000000 bcd_in2=00000110 cout=0 sum=00000110
* bcd_in1=00000000 bcd_in2=00000111 cout=0 sum=00000111
* bcd_in1=00000000 bcd_in2=00001000 cout=0 sum=00001000
* bcd_in1=00000000 bcd_in2=00001001 cout=0 sum=00001001
* bcd_in1=00000000 bcd_in2=00010000 cout=0 sum=00010000
* bcd_in1=00000000 bcd_in2=00010001 cout=0 sum=00010001
* bcd_in1=00000000 bcd_in2=00010010 cout=0 sum=00010010
* bcd_in1=00000000 bcd_in2=00010011 cout=0 sum=00010011
* bcd_in1=00000000 bcd_in2=00010100 cout=0 sum=00010100
* bcd_in1=00000000 bcd_in2=00010101 cout=0 sum=00010101
* bcd_in1=00000000 bcd_in2=00010110 cout=0 sum=00010110
* bcd_in1=00000000 bcd_in2=00010111 cout=0 sum=00010111
* bcd_in1=00000000 bcd_in2=00011000 cout=0 sum=00011000
* bcd_in1=00000000 bcd_in2=00011001 cout=0 sum=00011001
* bcd_in1=00000000 bcd_in2=00100000 cout=0 sum=00100000
* bcd_in1=00000000 bcd_in2=00100001 cout=0 sum=00100001
* bcd_in1=00000000 bcd_in2=00100010 cout=0 sum=00100010
* bcd_in1=00000000 bcd_in2=00100011 cout=0 sum=00100011
* bcd_in1=00000000 bcd_in2=00100100 cout=0 sum=00100100
* bcd_in1=00000000 bcd_in2=00100101 cout=0 sum=00100101
* bcd_in1=00000000 bcd_in2=00100110 cout=0 sum=00100110
* bcd_in1=00000000 bcd_in2=00100111 cout=0 sum=00100111
* bcd_in1=00000000 bcd_in2=00101000 cout=0 sum=00101000
* bcd_in1=00000000 bcd_in2=00101001 cout=0 sum=00101001
* bcd_in1=00000000 bcd_in2=00110000 cout=0 sum=00110000
* bcd_in1=00000000 bcd_in2=00110001 cout=0 sum=00110001
* bcd_in1=00000000 bcd_in2=00110010 cout=0 sum=00110010
* bcd_in1=00000000 bcd_in2=00110011 cout=0 sum=00110011
* bcd_in1=00000000 bcd_in2=00110100 cout=0 sum=00110100
* bcd_in1=00000000 bcd_in2=00110101 cout=0 sum=00110101
* bcd_in1=00000000 bcd_in2=00110110 cout=0 sum=00110110
* bcd_in1=00000000 bcd_in2=00110111 cout=0 sum=00110111
* bcd_in1=00000000 bcd_in2=00111000 cout=0 sum=00111000
* bcd_in1=00000000 bcd_in2=00111001 cout=0 sum=00111001
* bcd_in1=00000000 bcd_in2=01000000 cout=0 sum=01000000
* bcd_in1=00000000 bcd_in2=01000001 cout=0 sum=01000001
* bcd_in1=00000000 bcd_in2=01000010 cout=0 sum=01000010
* bcd_in1=00000000 bcd_in2=01000011 cout=0 sum=01000011
* bcd_in1=00000000 bcd_in2=01000100 cout=0 sum=01000100
* bcd_in1=00000000 bcd_in2=01000101 cout=0 sum=01000101
* bcd_in1=00000000 bcd_in2=01000110 cout=0 sum=01000110
* bcd_in1=00000000 bcd_in2=01000111 cout=0 sum=01000111
* bcd_in1=00000000 bcd_in2=01001000 cout=0 sum=01001000
* bcd_in1=00000000 bcd_in2=01001001 cout=0 sum=01001001
* bcd_in1=00000000 bcd_in2=01010000 cout=0 sum=01010000
* bcd_in1=00000000 bcd_in2=01010001 cout=0 sum=01010001
* bcd_in1=00000000 bcd_in2=01010010 cout=0 sum=01010010
* bcd_in1=00000000 bcd_in2=01010011 cout=0 sum=01010011
* bcd_in1=00000000 bcd_in2=01010100 cout=0 sum=01010100
* bcd_in1=00000000 bcd_in2=01010101 cout=0 sum=01010101
* bcd_in1=00000000 bcd_in2=01010110 cout=0 sum=01010110
* bcd_in1=00000000 bcd_in2=01010111 cout=0 sum=01010111
* bcd_in1=00000000 bcd_in2=01011000 cout=0 sum=01011000
* bcd_in1=00000000 bcd_in2=01011001 cout=0 sum=01011001
* bcd_in1=00000000 bcd_in2=01100000 cout=0 sum=01100000
* bcd_in1=00000000 bcd_in2=01100001 cout=0 sum=01100001
* bcd_in1=00000000 bcd_in2=01100010 cout=0 sum=01100010
* bcd_in1=00000000 bcd_in2=01100011 cout=0 sum=01100011
* bcd_in1=00000000 bcd_in2=01100100 cout=0 sum=01100100
* bcd_in1=00000000 bcd_in2=01100101 cout=0 sum=01100101
* bcd_in1=00000000 bcd_in2=01100110 cout=0 sum=01100110
* bcd_in1=00000000 bcd_in2=01100111 cout=0 sum=01100111
* bcd_in1=00000000 bcd_in2=01101000 cout=0 sum=01101000
* bcd_in1=00000000 bcd_in2=01101001 cout=0 sum=01101001
* bcd_in1=00000000 bcd_in2=01110000 cout=0 sum=01110000
* bcd_in1=00000000 bcd_in2=01110001 cout=0 sum=01110001
* bcd_in1=00000000 bcd_in2=01110010 cout=0 sum=01110010
* bcd_in1=00000000 bcd_in2=01110011 cout=0 sum=01110011
* bcd_in1=00000000 bcd_in2=01110100 cout=0 sum=01110100
* bcd_in1=00000000 bcd_in2=01110101 cout=0 sum=01110101
* bcd_in1=00000000 bcd_in2=01110110 cout=0 sum=01110110
* bcd_in1=00000000 bcd_in2=01110111 cout=0 sum=01110111
* bcd_in1=00000000 bcd_in2=01111000 cout=0 sum=01111000
* bcd_in1=00000000 bcd_in2=01111001 cout=0 sum=01111001
* bcd_in1=00000000 bcd_in2=10000000 cout=0 sum=10000000
* bcd_in1=00000000 bcd_in2=10000001 cout=0 sum=10000001
* bcd_in1=00000000 bcd_in2=10000010 cout=0 sum=10000010
* bcd_in1=00000000 bcd_in2=10000011 cout=0 sum=10000011
* bcd_in1=00000000 bcd_in2=10000100 cout=0 sum=10000100
* bcd_in1=00000000 bcd_in2=10000101 cout=0 sum=10000101
* bcd_in1=00000000 bcd_in2=10000110 cout=0 sum=10000110
* bcd_in1=00000000 bcd_in2=10000111 cout=0 sum=10000111
* bcd_in1=00000000 bcd_in2=10001000 cout=0 sum=10001000
* bcd_in1=00000000 bcd_in2=10001001 cout=0 sum=10001001
* bcd_in1=00000000 bcd_in2=10010000 cout=0 sum=10010000
* bcd_in1=00000000 bcd_in2=10010001 cout=0 sum=10010001
* bcd_in1=00000000 bcd_in2=10010010 cout=0 sum=10010010
* bcd_in1=00000000 bcd_in2=10010011 cout=0 sum=10010011
* bcd_in1=00000000 bcd_in2=10010100 cout=0 sum=10010100
* bcd_in1=00000000 bcd_in2=10010101 cout=0 sum=10010101
* bcd_in1=00000000 bcd_in2=10010110 cout=0 sum=10010110
* bcd_in1=00000000 bcd_in2=10010111 cout=0 sum=10010111
* bcd_in1=00000000 bcd_in2=10011000 cout=0 sum=10011000
* bcd_in1=00000000 bcd_in2=10011001 cout=0 sum=10011001
* bcd_in1=00000001 bcd_in2=00000000 cout=0 sum=00000001
* bcd_in1=00000001 bcd_in2=00000001 cout=0 sum=00000010
* bcd_in1=00000001 bcd_in2=00000010 cout=0 sum=00000011
* bcd_in1=00000001 bcd_in2=00000011 cout=0 sum=00000100
* bcd_in1=00000001 bcd_in2=00000100 cout=0 sum=00000101
* bcd_in1=00000001 bcd_in2=00000101 cout=0 sum=00000110
* bcd_in1=00000001 bcd_in2=00000110 cout=0 sum=00000111
* bcd_in1=00000001 bcd_in2=00000111 cout=0 sum=00001000
* bcd_in1=00000001 bcd_in2=00001000 cout=0 sum=00001001
* bcd_in1=00000001 bcd_in2=00001001 cout=0 sum=00010000
* bcd_in1=00000001 bcd_in2=00010000 cout=0 sum=00010001
* bcd_in1=00000001 bcd_in2=00010001 cout=0 sum=00010010
* bcd_in1=00000001 bcd_in2=00010010 cout=0 sum=00010011
* bcd_in1=00000001 bcd_in2=00010011 cout=0 sum=00010100
* bcd_in1=00000001 bcd_in2=00010100 cout=0 sum=00010101
* bcd_in1=00000001 bcd_in2=00010101 cout=0 sum=00010110
* bcd_in1=00000001 bcd_in2=00010110 cout=0 sum=00010111
* bcd_in1=00000001 bcd_in2=00010111 cout=0 sum=00011000
* bcd_in1=00000001 bcd_in2=00011000 cout=0 sum=00011001
* bcd_in1=00000001 bcd_in2=00011001 cout=0 sum=00100000
* bcd_in1=00000001 bcd_in2=00100000 cout=0 sum=00100001
* bcd_in1=00000001 bcd_in2=00100001 cout=0 sum=00100010
* bcd_in1=00000001 bcd_in2=00100010 cout=0 sum=00100011
* bcd_in1=00000001 bcd_in2=00100011 cout=0 sum=00100100
* bcd_in1=00000001 bcd_in2=00100100 cout=0 sum=00100101
* bcd_in1=00000001 bcd_in2=00100101 cout=0 sum=00100110
* bcd_in1=00000001 bcd_in2=00100110 cout=0 sum=00100111
* bcd_in1=00000001 bcd_in2=00100111 cout=0 sum=00101000
* bcd_in1=00000001 bcd_in2=00101000 cout=0 sum=00101001
* bcd_in1=00000001 bcd_in2=00101001 cout=0 sum=00110000
* bcd_in1=00000001 bcd_in2=00110000 cout=0 sum=00110001
* bcd_in1=00000001 bcd_in2=00110001 cout=0 sum=00110010
* bcd_in1=00000001 bcd_in2=00110010 cout=0 sum=00110011
* bcd_in1=00000001 bcd_in2=00110011 cout=0 sum=00110100
* bcd_in1=00000001 bcd_in2=00110100 cout=0 sum=00110101
* bcd_in1=00000001 bcd_in2=00110101 cout=0 sum=00110110
* bcd_in1=00000001 bcd_in2=00110110 cout=0 sum=00110111
* bcd_in1=00000001 bcd_in2=00110111 cout=0 sum=00111000
* bcd_in1=00000001 bcd_in2=00111000 cout=0 sum=00111001
* bcd_in1=00000001 bcd_in2=00111001 cout=0 sum=01000000
* bcd_in1=00000001 bcd_in2=01000000 cout=0 sum=01000001
* bcd_in1=00000001 bcd_in2=01000001 cout=0 sum=01000010
* bcd_in1=00000001 bcd_in2=01000010 cout=0 sum=01000011
* bcd_in1=00000001 bcd_in2=01000011 cout=0 sum=01000100
* bcd_in1=00000001 bcd_in2=01000100 cout=0 sum=01000101
* bcd_in1=00000001 bcd_in2=01000101 cout=0 sum=01000110
* bcd_in1=00000001 bcd_in2=01000110 cout=0 sum=01000111
* bcd_in1=00000001 bcd_in2=01000111 cout=0 sum=01001000
* bcd_in1=00000001 bcd_in2=01001000 cout=0 sum=01001001
* bcd_in1=00000001 bcd_in2=01001001 cout=0 sum=01010000
* bcd_in1=00000001 bcd_in2=01010000 cout=0 sum=01010001
* bcd_in1=00000001 bcd_in2=01010001 cout=0 sum=01010010
* bcd_in1=00000001 bcd_in2=01010010 cout=0 sum=01010011
* bcd_in1=00000001 bcd_in2=01010011 cout=0 sum=01010100
* bcd_in1=00000001 bcd_in2=01010100 cout=0 sum=01010101
* bcd_in1=00000001 bcd_in2=01010101 cout=0 sum=01010110
* bcd_in1=00000001 bcd_in2=01010110 cout=0 sum=01010111
* bcd_in1=00000001 bcd_in2=01010111 cout=0 sum=01011000
* bcd_in1=00000001 bcd_in2=01011000 cout=0 sum=01011001
* bcd_in1=00000001 bcd_in2=01011001 cout=0 sum=01100000
* bcd_in1=00000001 bcd_in2=01100000 cout=0 sum=01100001
* bcd_in1=00000001 bcd_in2=01100001 cout=0 sum=01100010
* bcd_in1=00000001 bcd_in2=01100010 cout=0 sum=01100011
* bcd_in1=00000001 bcd_in2=01100011 cout=0 sum=01100100
* bcd_in1=00000001 bcd_in2=01100100 cout=0 sum=01100101
* bcd_in1=00000001 bcd_in2=01100101 cout=0 sum=01100110
* bcd_in1=00000001 bcd_in2=01100110 cout=0 sum=01100111
* bcd_in1=00000001 bcd_in2=01100111 cout=0 sum=01101000
* bcd_in1=00000001 bcd_in2=01101000 cout=0 sum=01101001
* bcd_in1=00000001 bcd_in2=01101001 cout=0 sum=01110000
* bcd_in1=00000001 bcd_in2=01110000 cout=0 sum=01110001
* bcd_in1=00000001 bcd_in2=01110001 cout=0 sum=01110010
* bcd_in1=00000001 bcd_in2=01110010 cout=0 sum=01110011
* bcd_in1=00000001 bcd_in2=01110011 cout=0 sum=01110100
* bcd_in1=00000001 bcd_in2=01110100 cout=0 sum=01110101
* bcd_in1=00000001 bcd_in2=01110101 cout=0 sum=01110110
* bcd_in1=00000001 bcd_in2=01110110 cout=0 sum=01110111
* bcd_in1=00000001 bcd_in2=01110111 cout=0 sum=01111000
* bcd_in1=00000001 bcd_in2=01111000 cout=0 sum=01111001
* bcd_in1=00000001 bcd_in2=01111001 cout=0 sum=10000000
* bcd_in1=00000001 bcd_in2=10000000 cout=0 sum=10000001
* bcd_in1=00000001 bcd_in2=10000001 cout=0 sum=10000010
* bcd_in1=00000001 bcd_in2=10000010 cout=0 sum=10000011
* bcd_in1=00000001 bcd_in2=10000011 cout=0 sum=10000100
* bcd_in1=00000001 bcd_in2=10000100 cout=0 sum=10000101
* bcd_in1=00000001 bcd_in2=10000101 cout=0 sum=10000110
* bcd_in1=00000001 bcd_in2=10000110 cout=0 sum=10000111
* bcd_in1=00000001 bcd_in2=10000111 cout=0 sum=10001000
* bcd_in1=00000001 bcd_in2=10001000 cout=0 sum=10001001
* bcd_in1=00000001 bcd_in2=10001001 cout=0 sum=10010000
* bcd_in1=00000001 bcd_in2=10010000 cout=0 sum=10010001
* bcd_in1=00000001 bcd_in2=10010001 cout=0 sum=10010010
* bcd_in1=00000001 bcd_in2=10010010 cout=0 sum=10010011
* bcd_in1=00000001 bcd_in2=10010011 cout=0 sum=10010100
* bcd_in1=00000001 bcd_in2=10010100 cout=0 sum=10010101
* bcd_in1=00000001 bcd_in2=10010101 cout=0 sum=10010110
* bcd_in1=00000001 bcd_in2=10010110 cout=0 sum=10010111
* bcd_in1=00000001 bcd_in2=10010111 cout=0 sum=10011000
* bcd_in1=00000001 bcd_in2=10011000 cout=0 sum=10011001
* bcd_in1=00000001 bcd_in2=10011001 cout=1 sum=00000000
* bcd_in1=00000010 bcd_in2=00000000 cout=0 sum=00000010
* bcd_in1=00000010 bcd_in2=00000001 cout=0 sum=00000011
* bcd_in1=00000010 bcd_in2=00000010 cout=0 sum=00000100
* bcd_in1=00000010 bcd_in2=00000011 cout=0 sum=00000101
* bcd_in1=00000010 bcd_in2=00000100 cout=0 sum=00000110
* bcd_in1=00000010 bcd_in2=00000101 cout=0 sum=00000111
* bcd_in1=00000010 bcd_in2=00000110 cout=0 sum=00001000
* bcd_in1=00000010 bcd_in2=00000111 cout=0 sum=00001001
* bcd_in1=00000010 bcd_in2=00001000 cout=0 sum=00010000
* bcd_in1=00000010 bcd_in2=00001001 cout=0 sum=00010001
* bcd_in1=00000010 bcd_in2=00010000 cout=0 sum=00010010
* bcd_in1=00000010 bcd_in2=00010001 cout=0 sum=00010011
* bcd_in1=00000010 bcd_in2=00010010 cout=0 sum=00010100
* bcd_in1=00000010 bcd_in2=00010011 cout=0 sum=00010101
* bcd_in1=00000010 bcd_in2=00010100 cout=0 sum=00010110
* bcd_in1=00000010 bcd_in2=00010101 cout=0 sum=00010111
* bcd_in1=00000010 bcd_in2=00010110 cout=0 sum=00011000
* bcd_in1=00000010 bcd_in2=00010111 cout=0 sum=00011001
* bcd_in1=00000010 bcd_in2=00011000 cout=0 sum=00100000
* bcd_in1=00000010 bcd_in2=00011001 cout=0 sum=00100001
* bcd_in1=00000010 bcd_in2=00100000 cout=0 sum=00100010
* bcd_in1=00000010 bcd_in2=00100001 cout=0 sum=00100011
* bcd_in1=00000010 bcd_in2=00100010 cout=0 sum=00100100
* bcd_in1=00000010 bcd_in2=00100011 cout=0 sum=00100101
* bcd_in1=00000010 bcd_in2=00100100 cout=0 sum=00100110
* bcd_in1=00000010 bcd_in2=00100101 cout=0 sum=00100111
* bcd_in1=00000010 bcd_in2=00100110 cout=0 sum=00101000
* bcd_in1=00000010 bcd_in2=00100111 cout=0 sum=00101001
* bcd_in1=00000010 bcd_in2=00101000 cout=0 sum=00110000
* bcd_in1=00000010 bcd_in2=00101001 cout=0 sum=00110001
* bcd_in1=00000010 bcd_in2=00110000 cout=0 sum=00110010
* bcd_in1=00000010 bcd_in2=00110001 cout=0 sum=00110011
* bcd_in1=00000010 bcd_in2=00110010 cout=0 sum=00110100
* bcd_in1=00000010 bcd_in2=00110011 cout=0 sum=00110101
* bcd_in1=00000010 bcd_in2=00110100 cout=0 sum=00110110
* bcd_in1=00000010 bcd_in2=00110101 cout=0 sum=00110111
* bcd_in1=00000010 bcd_in2=00110110 cout=0 sum=00111000
* bcd_in1=00000010 bcd_in2=00110111 cout=0 sum=00111001
* bcd_in1=00000010 bcd_in2=00111000 cout=0 sum=01000000
* bcd_in1=00000010 bcd_in2=00111001 cout=0 sum=01000001
* bcd_in1=00000010 bcd_in2=01000000 cout=0 sum=01000010
* bcd_in1=00000010 bcd_in2=01000001 cout=0 sum=01000011
* bcd_in1=00000010 bcd_in2=01000010 cout=0 sum=01000100
* bcd_in1=00000010 bcd_in2=01000011 cout=0 sum=01000101
* bcd_in1=00000010 bcd_in2=01000100 cout=0 sum=01000110
* bcd_in1=00000010 bcd_in2=01000101 cout=0 sum=01000111
* bcd_in1=00000010 bcd_in2=01000110 cout=0 sum=01001000
* bcd_in1=00000010 bcd_in2=01000111 cout=0 sum=01001001
* bcd_in1=00000010 bcd_in2=01001000 cout=0 sum=01010000
* bcd_in1=00000010 bcd_in2=01001001 cout=0 sum=01010001
* bcd_in1=00000010 bcd_in2=01010000 cout=0 sum=01010010
* bcd_in1=00000010 bcd_in2=01010001 cout=0 sum=01010011
* bcd_in1=00000010 bcd_in2=01010010 cout=0 sum=01010100
* bcd_in1=00000010 bcd_in2=01010011 cout=0 sum=01010101
* bcd_in1=00000010 bcd_in2=01010100 cout=0 sum=01010110
* bcd_in1=00000010 bcd_in2=01010101 cout=0 sum=01010111
* bcd_in1=00000010 bcd_in2=01010110 cout=0 sum=01011000
* bcd_in1=00000010 bcd_in2=01010111 cout=0 sum=01011001
* bcd_in1=00000010 bcd_in2=01011000 cout=0 sum=01100000
* bcd_in1=00000010 bcd_in2=01011001 cout=0 sum=01100001
* bcd_in1=00000010 bcd_in2=01100000 cout=0 sum=01100010
* bcd_in1=00000010 bcd_in2=01100001 cout=0 sum=01100011
* bcd_in1=00000010 bcd_in2=01100010 cout=0 sum=01100100
* bcd_in1=00000010 bcd_in2=01100011 cout=0 sum=01100101
* bcd_in1=00000010 bcd_in2=01100100 cout=0 sum=01100110
* bcd_in1=00000010 bcd_in2=01100101 cout=0 sum=01100111
* bcd_in1=00000010 bcd_in2=01100110 cout=0 sum=01101000
* bcd_in1=00000010 bcd_in2=01100111 cout=0 sum=01101001
* bcd_in1=00000010 bcd_in2=01101000 cout=0 sum=01110000
* bcd_in1=00000010 bcd_in2=01101001 cout=0 sum=01110001
* bcd_in1=00000010 bcd_in2=01110000 cout=0 sum=01110010
* bcd_in1=00000010 bcd_in2=01110001 cout=0 sum=01110011
* bcd_in1=00000010 bcd_in2=01110010 cout=0 sum=01110100
* bcd_in1=00000010 bcd_in2=01110011 cout=0 sum=01110101
* bcd_in1=00000010 bcd_in2=01110100 cout=0 sum=01110110
* bcd_in1=00000010 bcd_in2=01110101 cout=0 sum=01110111
* bcd_in1=00000010 bcd_in2=01110110 cout=0 sum=01111000
* bcd_in1=00000010 bcd_in2=01110111 cout=0 sum=01111001
* bcd_in1=00000010 bcd_in2=01111000 cout=0 sum=10000000
* bcd_in1=00000010 bcd_in2=01111001 cout=0 sum=10000001
* bcd_in1=00000010 bcd_in2=10000000 cout=0 sum=10000010
* bcd_in1=00000010 bcd_in2=10000001 cout=0 sum=10000011
* bcd_in1=00000010 bcd_in2=10000010 cout=0 sum=10000100
* bcd_in1=00000010 bcd_in2=10000011 cout=0 sum=10000101
* bcd_in1=00000010 bcd_in2=10000100 cout=0 sum=10000110
* bcd_in1=00000010 bcd_in2=10000101 cout=0 sum=10000111
* bcd_in1=00000010 bcd_in2=10000110 cout=0 sum=10001000
* bcd_in1=00000010 bcd_in2=10000111 cout=0 sum=10001001
* bcd_in1=00000010 bcd_in2=10001000 cout=0 sum=10010000
* bcd_in1=00000010 bcd_in2=10001001 cout=0 sum=10010001
* bcd_in1=00000010 bcd_in2=10010000 cout=0 sum=10010010
* bcd_in1=00000010 bcd_in2=10010001 cout=0 sum=10010011
* bcd_in1=00000010 bcd_in2=10010010 cout=0 sum=10010100
* bcd_in1=00000010 bcd_in2=10010011 cout=0 sum=10010101
* bcd_in1=00000010 bcd_in2=10010100 cout=0 sum=10010110
* bcd_in1=00000010 bcd_in2=10010101 cout=0 sum=10010111
* bcd_in1=00000010 bcd_in2=10010110 cout=0 sum=10011000
* bcd_in1=00000010 bcd_in2=10010111 cout=0 sum=10011001
* bcd_in1=00000010 bcd_in2=10011000 cout=1 sum=00000000
* bcd_in1=00000010 bcd_in2=10011001 cout=1 sum=00000001
* bcd_in1=00000011 bcd_in2=00000000 cout=0 sum=00000011
* bcd_in1=00000011 bcd_in2=00000001 cout=0 sum=00000100
* bcd_in1=00000011 bcd_in2=00000010 cout=0 sum=00000101
* bcd_in1=00000011 bcd_in2=00000011 cout=0 sum=00000110
* bcd_in1=00000011 bcd_in2=00000100 cout=0 sum=00000111
* bcd_in1=00000011 bcd_in2=00000101 cout=0 sum=00001000
* bcd_in1=00000011 bcd_in2=00000110 cout=0 sum=00001001
* bcd_in1=00000011 bcd_in2=00000111 cout=0 sum=00010000
* bcd_in1=00000011 bcd_in2=00001000 cout=0 sum=00010001
* bcd_in1=00000011 bcd_in2=00001001 cout=0 sum=00010010
* bcd_in1=00000011 bcd_in2=00010000 cout=0 sum=00010011
* bcd_in1=00000011 bcd_in2=00010001 cout=0 sum=00010100
* bcd_in1=00000011 bcd_in2=00010010 cout=0 sum=00010101
* bcd_in1=00000011 bcd_in2=00010011 cout=0 sum=00010110
* bcd_in1=00000011 bcd_in2=00010100 cout=0 sum=00010111
* bcd_in1=00000011 bcd_in2=00010101 cout=0 sum=00011000
* bcd_in1=00000011 bcd_in2=00010110 cout=0 sum=00011001
* bcd_in1=00000011 bcd_in2=00010111 cout=0 sum=00100000
* bcd_in1=00000011 bcd_in2=00011000 cout=0 sum=00100001
* bcd_in1=00000011 bcd_in2=00011001 cout=0 sum=00100010
* bcd_in1=00000011 bcd_in2=00100000 cout=0 sum=00100011
* bcd_in1=00000011 bcd_in2=00100001 cout=0 sum=00100100
* bcd_in1=00000011 bcd_in2=00100010 cout=0 sum=00100101
* bcd_in1=00000011 bcd_in2=00100011 cout=0 sum=00100110
* bcd_in1=00000011 bcd_in2=00100100 cout=0 sum=00100111
* bcd_in1=00000011 bcd_in2=00100101 cout=0 sum=00101000
* bcd_in1=00000011 bcd_in2=00100110 cout=0 sum=00101001
* bcd_in1=00000011 bcd_in2=00100111 cout=0 sum=00110000
* bcd_in1=00000011 bcd_in2=00101000 cout=0 sum=00110001
* bcd_in1=00000011 bcd_in2=00101001 cout=0 sum=00110010
* bcd_in1=00000011 bcd_in2=00110000 cout=0 sum=00110011
* bcd_in1=00000011 bcd_in2=00110001 cout=0 sum=00110100
* bcd_in1=00000011 bcd_in2=00110010 cout=0 sum=00110101
* bcd_in1=00000011 bcd_in2=00110011 cout=0 sum=00110110
* bcd_in1=00000011 bcd_in2=00110100 cout=0 sum=00110111
* bcd_in1=00000011 bcd_in2=00110101 cout=0 sum=00111000
* bcd_in1=00000011 bcd_in2=00110110 cout=0 sum=00111001
* bcd_in1=00000011 bcd_in2=00110111 cout=0 sum=01000000
* bcd_in1=00000011 bcd_in2=00111000 cout=0 sum=01000001
* bcd_in1=00000011 bcd_in2=00111001 cout=0 sum=01000010
* bcd_in1=00000011 bcd_in2=01000000 cout=0 sum=01000011
* bcd_in1=00000011 bcd_in2=01000001 cout=0 sum=01000100
* bcd_in1=00000011 bcd_in2=01000010 cout=0 sum=01000101
* bcd_in1=00000011 bcd_in2=01000011 cout=0 sum=01000110
* bcd_in1=00000011 bcd_in2=01000100 cout=0 sum=01000111
* bcd_in1=00000011 bcd_in2=01000101 cout=0 sum=01001000
* bcd_in1=00000011 bcd_in2=01000110 cout=0 sum=01001001
* bcd_in1=00000011 bcd_in2=01000111 cout=0 sum=01010000
* bcd_in1=00000011 bcd_in2=01001000 cout=0 sum=01010001
* bcd_in1=00000011 bcd_in2=01001001 cout=0 sum=01010010
* bcd_in1=00000011 bcd_in2=01010000 cout=0 sum=01010011
* bcd_in1=00000011 bcd_in2=01010001 cout=0 sum=01010100
* bcd_in1=00000011 bcd_in2=01010010 cout=0 sum=01010101
* bcd_in1=00000011 bcd_in2=01010011 cout=0 sum=01010110
* bcd_in1=00000011 bcd_in2=01010100 cout=0 sum=01010111
* bcd_in1=00000011 bcd_in2=01010101 cout=0 sum=01011000
* bcd_in1=00000011 bcd_in2=01010110 cout=0 sum=01011001
* bcd_in1=00000011 bcd_in2=01010111 cout=0 sum=01100000
* bcd_in1=00000011 bcd_in2=01011000 cout=0 sum=01100001
* bcd_in1=00000011 bcd_in2=01011001 cout=0 sum=01100010
* bcd_in1=00000011 bcd_in2=01100000 cout=0 sum=01100011
* bcd_in1=00000011 bcd_in2=01100001 cout=0 sum=01100100
* bcd_in1=00000011 bcd_in2=01100010 cout=0 sum=01100101
* bcd_in1=00000011 bcd_in2=01100011 cout=0 sum=01100110
* bcd_in1=00000011 bcd_in2=01100100 cout=0 sum=01100111
* bcd_in1=00000011 bcd_in2=01100101 cout=0 sum=01101000
* bcd_in1=00000011 bcd_in2=01100110 cout=0 sum=01101001
* bcd_in1=00000011 bcd_in2=01100111 cout=0 sum=01110000
* bcd_in1=00000011 bcd_in2=01101000 cout=0 sum=01110001
* bcd_in1=00000011 bcd_in2=01101001 cout=0 sum=01110010
* bcd_in1=00000011 bcd_in2=01110000 cout=0 sum=01110011
* bcd_in1=00000011 bcd_in2=01110001 cout=0 sum=01110100
* bcd_in1=00000011 bcd_in2=01110010 cout=0 sum=01110101
* bcd_in1=00000011 bcd_in2=01110011 cout=0 sum=01110110
* bcd_in1=00000011 bcd_in2=01110100 cout=0 sum=01110111
* bcd_in1=00000011 bcd_in2=01110101 cout=0 sum=01111000
* bcd_in1=00000011 bcd_in2=01110110 cout=0 sum=01111001
* bcd_in1=00000011 bcd_in2=01110111 cout=0 sum=10000000
* bcd_in1=00000011 bcd_in2=01111000 cout=0 sum=10000001
* bcd_in1=00000011 bcd_in2=01111001 cout=0 sum=10000010
* bcd_in1=00000011 bcd_in2=10000000 cout=0 sum=10000011
* bcd_in1=00000011 bcd_in2=10000001 cout=0 sum=10000100
* bcd_in1=00000011 bcd_in2=10000010 cout=0 sum=10000101
* bcd_in1=00000011 bcd_in2=10000011 cout=0 sum=10000110
* bcd_in1=00000011 bcd_in2=10000100 cout=0 sum=10000111
* bcd_in1=00000011 bcd_in2=10000101 cout=0 sum=10001000
* bcd_in1=00000011 bcd_in2=10000110 cout=0 sum=10001001
* bcd_in1=00000011 bcd_in2=10000111 cout=0 sum=10010000
* bcd_in1=00000011 bcd_in2=10001000 cout=0 sum=10010001
* bcd_in1=00000011 bcd_in2=10001001 cout=0 sum=10010010
* bcd_in1=00000011 bcd_in2=10010000 cout=0 sum=10010011
* bcd_in1=00000011 bcd_in2=10010001 cout=0 sum=10010100
* bcd_in1=00000011 bcd_in2=10010010 cout=0 sum=10010101
* bcd_in1=00000011 bcd_in2=10010011 cout=0 sum=10010110
* bcd_in1=00000011 bcd_in2=10010100 cout=0 sum=10010111
* bcd_in1=00000011 bcd_in2=10010101 cout=0 sum=10011000
* bcd_in1=00000011 bcd_in2=10010110 cout=0 sum=10011001
* bcd_in1=00000011 bcd_in2=10010111 cout=1 sum=00000000
* bcd_in1=00000011 bcd_in2=10011000 cout=1 sum=00000001
* bcd_in1=00000011 bcd_in2=10011001 cout=1 sum=00000010
* bcd_in1=00000100 bcd_in2=00000000 cout=0 sum=00000100
* bcd_in1=00000100 bcd_in2=00000001 cout=0 sum=00000101
* bcd_in1=00000100 bcd_in2=00000010 cout=0 sum=00000110
* bcd_in1=00000100 bcd_in2=00000011 cout=0 sum=00000111
* bcd_in1=00000100 bcd_in2=00000100 cout=0 sum=00001000
* bcd_in1=00000100 bcd_in2=00000101 cout=0 sum=00001001
* bcd_in1=00000100 bcd_in2=00000110 cout=0 sum=00010000
* bcd_in1=00000100 bcd_in2=00000111 cout=0 sum=00010001
* bcd_in1=00000100 bcd_in2=00001000 cout=0 sum=00010010
* bcd_in1=00000100 bcd_in2=00001001 cout=0 sum=00010011
* bcd_in1=00000100 bcd_in2=00010000 cout=0 sum=00010100
* bcd_in1=00000100 bcd_in2=00010001 cout=0 sum=00010101
* bcd_in1=00000100 bcd_in2=00010010 cout=0 sum=00010110
* bcd_in1=00000100 bcd_in2=00010011 cout=0 sum=00010111
* bcd_in1=00000100 bcd_in2=00010100 cout=0 sum=00011000
* bcd_in1=00000100 bcd_in2=00010101 cout=0 sum=00011001
* bcd_in1=00000100 bcd_in2=00010110 cout=0 sum=00100000
* bcd_in1=00000100 bcd_in2=00010111 cout=0 sum=00100001
* bcd_in1=00000100 bcd_in2=00011000 cout=0 sum=00100010
* bcd_in1=00000100 bcd_in2=00011001 cout=0 sum=00100011
* bcd_in1=00000100 bcd_in2=00100000 cout=0 sum=00100100
* bcd_in1=00000100 bcd_in2=00100001 cout=0 sum=00100101
* bcd_in1=00000100 bcd_in2=00100010 cout=0 sum=00100110
* bcd_in1=00000100 bcd_in2=00100011 cout=0 sum=00100111
* bcd_in1=00000100 bcd_in2=00100100 cout=0 sum=00101000
* bcd_in1=00000100 bcd_in2=00100101 cout=0 sum=00101001
* bcd_in1=00000100 bcd_in2=00100110 cout=0 sum=00110000
* bcd_in1=00000100 bcd_in2=00100111 cout=0 sum=00110001
* bcd_in1=00000100 bcd_in2=00101000 cout=0 sum=00110010
* bcd_in1=00000100 bcd_in2=00101001 cout=0 sum=00110011
* bcd_in1=00000100 bcd_in2=00110000 cout=0 sum=00110100
* bcd_in1=00000100 bcd_in2=00110001 cout=0 sum=00110101
* bcd_in1=00000100 bcd_in2=00110010 cout=0 sum=00110110
* bcd_in1=00000100 bcd_in2=00110011 cout=0 sum=00110111
* bcd_in1=00000100 bcd_in2=00110100 cout=0 sum=00111000
* bcd_in1=00000100 bcd_in2=00110101 cout=0 sum=00111001
* bcd_in1=00000100 bcd_in2=00110110 cout=0 sum=01000000
* bcd_in1=00000100 bcd_in2=00110111 cout=0 sum=01000001
* bcd_in1=00000100 bcd_in2=00111000 cout=0 sum=01000010
* bcd_in1=00000100 bcd_in2=00111001 cout=0 sum=01000011
* bcd_in1=00000100 bcd_in2=01000000 cout=0 sum=01000100
* bcd_in1=00000100 bcd_in2=01000001 cout=0 sum=01000101
* bcd_in1=00000100 bcd_in2=01000010 cout=0 sum=01000110
* bcd_in1=00000100 bcd_in2=01000011 cout=0 sum=01000111
* bcd_in1=00000100 bcd_in2=01000100 cout=0 sum=01001000
* bcd_in1=00000100 bcd_in2=01000101 cout=0 sum=01001001
* bcd_in1=00000100 bcd_in2=01000110 cout=0 sum=01010000
* bcd_in1=00000100 bcd_in2=01000111 cout=0 sum=01010001
* bcd_in1=00000100 bcd_in2=01001000 cout=0 sum=01010010
* bcd_in1=00000100 bcd_in2=01001001 cout=0 sum=01010011
* bcd_in1=00000100 bcd_in2=01010000 cout=0 sum=01010100
* bcd_in1=00000100 bcd_in2=01010001 cout=0 sum=01010101
* bcd_in1=00000100 bcd_in2=01010010 cout=0 sum=01010110
* bcd_in1=00000100 bcd_in2=01010011 cout=0 sum=01010111
* bcd_in1=00000100 bcd_in2=01010100 cout=0 sum=01011000
* bcd_in1=00000100 bcd_in2=01010101 cout=0 sum=01011001
* bcd_in1=00000100 bcd_in2=01010110 cout=0 sum=01100000
* bcd_in1=00000100 bcd_in2=01010111 cout=0 sum=01100001
* bcd_in1=00000100 bcd_in2=01011000 cout=0 sum=01100010
* bcd_in1=00000100 bcd_in2=01011001 cout=0 sum=01100011
* bcd_in1=00000100 bcd_in2=01100000 cout=0 sum=01100100
* bcd_in1=00000100 bcd_in2=01100001 cout=0 sum=01100101
* bcd_in1=00000100 bcd_in2=01100010 cout=0 sum=01100110
* bcd_in1=00000100 bcd_in2=01100011 cout=0 sum=01100111
* bcd_in1=00000100 bcd_in2=01100100 cout=0 sum=01101000
* bcd_in1=00000100 bcd_in2=01100101 cout=0 sum=01101001
* bcd_in1=00000100 bcd_in2=01100110 cout=0 sum=01110000
* bcd_in1=00000100 bcd_in2=01100111 cout=0 sum=01110001
* bcd_in1=00000100 bcd_in2=01101000 cout=0 sum=01110010
* bcd_in1=00000100 bcd_in2=01101001 cout=0 sum=01110011
* bcd_in1=00000100 bcd_in2=01110000 cout=0 sum=01110100
* bcd_in1=00000100 bcd_in2=01110001 cout=0 sum=01110101
* bcd_in1=00000100 bcd_in2=01110010 cout=0 sum=01110110
* bcd_in1=00000100 bcd_in2=01110011 cout=0 sum=01110111
* bcd_in1=00000100 bcd_in2=01110100 cout=0 sum=01111000
* bcd_in1=00000100 bcd_in2=01110101 cout=0 sum=01111001
* bcd_in1=00000100 bcd_in2=01110110 cout=0 sum=10000000
* bcd_in1=00000100 bcd_in2=01110111 cout=0 sum=10000001
* bcd_in1=00000100 bcd_in2=01111000 cout=0 sum=10000010
* bcd_in1=00000100 bcd_in2=01111001 cout=0 sum=10000011
* bcd_in1=00000100 bcd_in2=10000000 cout=0 sum=10000100
* bcd_in1=00000100 bcd_in2=10000001 cout=0 sum=10000101
* bcd_in1=00000100 bcd_in2=10000010 cout=0 sum=10000110
* bcd_in1=00000100 bcd_in2=10000011 cout=0 sum=10000111
* bcd_in1=00000100 bcd_in2=10000100 cout=0 sum=10001000
* bcd_in1=00000100 bcd_in2=10000101 cout=0 sum=10001001
* bcd_in1=00000100 bcd_in2=10000110 cout=0 sum=10010000
* bcd_in1=00000100 bcd_in2=10000111 cout=0 sum=10010001
* bcd_in1=00000100 bcd_in2=10001000 cout=0 sum=10010010
* bcd_in1=00000100 bcd_in2=10001001 cout=0 sum=10010011
* bcd_in1=00000100 bcd_in2=10010000 cout=0 sum=10010100
* bcd_in1=00000100 bcd_in2=10010001 cout=0 sum=10010101
* bcd_in1=00000100 bcd_in2=10010010 cout=0 sum=10010110
* bcd_in1=00000100 bcd_in2=10010011 cout=0 sum=10010111
* bcd_in1=00000100 bcd_in2=10010100 cout=0 sum=10011000
* bcd_in1=00000100 bcd_in2=10010101 cout=0 sum=10011001
* bcd_in1=00000100 bcd_in2=10010110 cout=1 sum=00000000
* bcd_in1=00000100 bcd_in2=10010111 cout=1 sum=00000001
* bcd_in1=00000100 bcd_in2=10011000 cout=1 sum=00000010
* bcd_in1=00000100 bcd_in2=10011001 cout=1 sum=00000011
* bcd_in1=00000101 bcd_in2=00000000 cout=0 sum=00000101
* bcd_in1=00000101 bcd_in2=00000001 cout=0 sum=00000110
* bcd_in1=00000101 bcd_in2=00000010 cout=0 sum=00000111
* bcd_in1=00000101 bcd_in2=00000011 cout=0 sum=00001000
* bcd_in1=00000101 bcd_in2=00000100 cout=0 sum=00001001
* bcd_in1=00000101 bcd_in2=00000101 cout=0 sum=00010000
* bcd_in1=00000101 bcd_in2=00000110 cout=0 sum=00010001
* bcd_in1=00000101 bcd_in2=00000111 cout=0 sum=00010010
* bcd_in1=00000101 bcd_in2=00001000 cout=0 sum=00010011
* bcd_in1=00000101 bcd_in2=00001001 cout=0 sum=00010100
* bcd_in1=00000101 bcd_in2=00010000 cout=0 sum=00010101
* bcd_in1=00000101 bcd_in2=00010001 cout=0 sum=00010110
* bcd_in1=00000101 bcd_in2=00010010 cout=0 sum=00010111
* bcd_in1=00000101 bcd_in2=00010011 cout=0 sum=00011000
* bcd_in1=00000101 bcd_in2=00010100 cout=0 sum=00011001
* bcd_in1=00000101 bcd_in2=00010101 cout=0 sum=00100000
* bcd_in1=00000101 bcd_in2=00010110 cout=0 sum=00100001
* bcd_in1=00000101 bcd_in2=00010111 cout=0 sum=00100010
* bcd_in1=00000101 bcd_in2=00011000 cout=0 sum=00100011
* bcd_in1=00000101 bcd_in2=00011001 cout=0 sum=00100100
* bcd_in1=00000101 bcd_in2=00100000 cout=0 sum=00100101
* bcd_in1=00000101 bcd_in2=00100001 cout=0 sum=00100110
* bcd_in1=00000101 bcd_in2=00100010 cout=0 sum=00100111
* bcd_in1=00000101 bcd_in2=00100011 cout=0 sum=00101000
* bcd_in1=00000101 bcd_in2=00100100 cout=0 sum=00101001
* bcd_in1=00000101 bcd_in2=00100101 cout=0 sum=00110000
* bcd_in1=00000101 bcd_in2=00100110 cout=0 sum=00110001
* bcd_in1=00000101 bcd_in2=00100111 cout=0 sum=00110010
* bcd_in1=00000101 bcd_in2=00101000 cout=0 sum=00110011
* bcd_in1=00000101 bcd_in2=00101001 cout=0 sum=00110100
* bcd_in1=00000101 bcd_in2=00110000 cout=0 sum=00110101
* bcd_in1=00000101 bcd_in2=00110001 cout=0 sum=00110110
* bcd_in1=00000101 bcd_in2=00110010 cout=0 sum=00110111
* bcd_in1=00000101 bcd_in2=00110011 cout=0 sum=00111000
* bcd_in1=00000101 bcd_in2=00110100 cout=0 sum=00111001
* bcd_in1=00000101 bcd_in2=00110101 cout=0 sum=01000000
* bcd_in1=00000101 bcd_in2=00110110 cout=0 sum=01000001
* bcd_in1=00000101 bcd_in2=00110111 cout=0 sum=01000010
* bcd_in1=00000101 bcd_in2=00111000 cout=0 sum=01000011
* bcd_in1=00000101 bcd_in2=00111001 cout=0 sum=01000100
* bcd_in1=00000101 bcd_in2=01000000 cout=0 sum=01000101
* bcd_in1=00000101 bcd_in2=01000001 cout=0 sum=01000110
* bcd_in1=00000101 bcd_in2=01000010 cout=0 sum=01000111
* bcd_in1=00000101 bcd_in2=01000011 cout=0 sum=01001000
* bcd_in1=00000101 bcd_in2=01000100 cout=0 sum=01001001
* bcd_in1=00000101 bcd_in2=01000101 cout=0 sum=01010000
* bcd_in1=00000101 bcd_in2=01000110 cout=0 sum=01010001
* bcd_in1=00000101 bcd_in2=01000111 cout=0 sum=01010010
* bcd_in1=00000101 bcd_in2=01001000 cout=0 sum=01010011
* bcd_in1=00000101 bcd_in2=01001001 cout=0 sum=01010100
* bcd_in1=00000101 bcd_in2=01010000 cout=0 sum=01010101
* bcd_in1=00000101 bcd_in2=01010001 cout=0 sum=01010110
* bcd_in1=00000101 bcd_in2=01010010 cout=0 sum=01010111
* bcd_in1=00000101 bcd_in2=01010011 cout=0 sum=01011000
* bcd_in1=00000101 bcd_in2=01010100 cout=0 sum=01011001
* bcd_in1=00000101 bcd_in2=01010101 cout=0 sum=01100000
* bcd_in1=00000101 bcd_in2=01010110 cout=0 sum=01100001
* bcd_in1=00000101 bcd_in2=01010111 cout=0 sum=01100010
* bcd_in1=00000101 bcd_in2=01011000 cout=0 sum=01100011
* bcd_in1=00000101 bcd_in2=01011001 cout=0 sum=01100100
* bcd_in1=00000101 bcd_in2=01100000 cout=0 sum=01100101
* bcd_in1=00000101 bcd_in2=01100001 cout=0 sum=01100110
* bcd_in1=00000101 bcd_in2=01100010 cout=0 sum=01100111
* bcd_in1=00000101 bcd_in2=01100011 cout=0 sum=01101000
* bcd_in1=00000101 bcd_in2=01100100 cout=0 sum=01101001
* bcd_in1=00000101 bcd_in2=01100101 cout=0 sum=01110000
* bcd_in1=00000101 bcd_in2=01100110 cout=0 sum=01110001
* bcd_in1=00000101 bcd_in2=01100111 cout=0 sum=01110010
* bcd_in1=00000101 bcd_in2=01101000 cout=0 sum=01110011
* bcd_in1=00000101 bcd_in2=01101001 cout=0 sum=01110100
* bcd_in1=00000101 bcd_in2=01110000 cout=0 sum=01110101
* bcd_in1=00000101 bcd_in2=01110001 cout=0 sum=01110110
* bcd_in1=00000101 bcd_in2=01110010 cout=0 sum=01110111
* bcd_in1=00000101 bcd_in2=01110011 cout=0 sum=01111000
* bcd_in1=00000101 bcd_in2=01110100 cout=0 sum=01111001
* bcd_in1=00000101 bcd_in2=01110101 cout=0 sum=10000000
* bcd_in1=00000101 bcd_in2=01110110 cout=0 sum=10000001
* bcd_in1=00000101 bcd_in2=01110111 cout=0 sum=10000010
* bcd_in1=00000101 bcd_in2=01111000 cout=0 sum=10000011
* bcd_in1=00000101 bcd_in2=01111001 cout=0 sum=10000100
* bcd_in1=00000101 bcd_in2=10000000 cout=0 sum=10000101
* bcd_in1=00000101 bcd_in2=10000001 cout=0 sum=10000110
* bcd_in1=00000101 bcd_in2=10000010 cout=0 sum=10000111
* bcd_in1=00000101 bcd_in2=10000011 cout=0 sum=10001000
* bcd_in1=00000101 bcd_in2=10000100 cout=0 sum=10001001
* bcd_in1=00000101 bcd_in2=10000101 cout=0 sum=10010000
* bcd_in1=00000101 bcd_in2=10000110 cout=0 sum=10010001
* bcd_in1=00000101 bcd_in2=10000111 cout=0 sum=10010010
* bcd_in1=00000101 bcd_in2=10001000 cout=0 sum=10010011
* bcd_in1=00000101 bcd_in2=10001001 cout=0 sum=10010100
* bcd_in1=00000101 bcd_in2=10010000 cout=0 sum=10010101
* bcd_in1=00000101 bcd_in2=10010001 cout=0 sum=10010110
* bcd_in1=00000101 bcd_in2=10010010 cout=0 sum=10010111
* bcd_in1=00000101 bcd_in2=10010011 cout=0 sum=10011000
* bcd_in1=00000101 bcd_in2=10010100 cout=0 sum=10011001
* bcd_in1=00000101 bcd_in2=10010101 cout=1 sum=00000000
* bcd_in1=00000101 bcd_in2=10010110 cout=1 sum=00000001
* bcd_in1=00000101 bcd_in2=10010111 cout=1 sum=00000010
* bcd_in1=00000101 bcd_in2=10011000 cout=1 sum=00000011
* bcd_in1=00000101 bcd_in2=10011001 cout=1 sum=00000100
* bcd_in1=00000110 bcd_in2=00000000 cout=0 sum=00000110
* bcd_in1=00000110 bcd_in2=00000001 cout=0 sum=00000111
* bcd_in1=00000110 bcd_in2=00000010 cout=0 sum=00001000
* bcd_in1=00000110 bcd_in2=00000011 cout=0 sum=00001001
* bcd_in1=00000110 bcd_in2=00000100 cout=0 sum=00010000
* bcd_in1=00000110 bcd_in2=00000101 cout=0 sum=00010001
* bcd_in1=00000110 bcd_in2=00000110 cout=0 sum=00010010
* bcd_in1=00000110 bcd_in2=00000111 cout=0 sum=00010011
* bcd_in1=00000110 bcd_in2=00001000 cout=0 sum=00010100
* bcd_in1=00000110 bcd_in2=00001001 cout=0 sum=00010101
* bcd_in1=00000110 bcd_in2=00010000 cout=0 sum=00010110
* bcd_in1=00000110 bcd_in2=00010001 cout=0 sum=00010111
* bcd_in1=00000110 bcd_in2=00010010 cout=0 sum=00011000
* bcd_in1=00000110 bcd_in2=00010011 cout=0 sum=00011001
* bcd_in1=00000110 bcd_in2=00010100 cout=0 sum=00100000
* bcd_in1=00000110 bcd_in2=00010101 cout=0 sum=00100001
* bcd_in1=00000110 bcd_in2=00010110 cout=0 sum=00100010
* bcd_in1=00000110 bcd_in2=00010111 cout=0 sum=00100011
* bcd_in1=00000110 bcd_in2=00011000 cout=0 sum=00100100
* bcd_in1=00000110 bcd_in2=00011001 cout=0 sum=00100101
* bcd_in1=00000110 bcd_in2=00100000 cout=0 sum=00100110
* bcd_in1=00000110 bcd_in2=00100001 cout=0 sum=00100111
* bcd_in1=00000110 bcd_in2=00100010 cout=0 sum=00101000
* bcd_in1=00000110 bcd_in2=00100011 cout=0 sum=00101001
* bcd_in1=00000110 bcd_in2=00100100 cout=0 sum=00110000
* bcd_in1=00000110 bcd_in2=00100101 cout=0 sum=00110001
* bcd_in1=00000110 bcd_in2=00100110 cout=0 sum=00110010
* bcd_in1=00000110 bcd_in2=00100111 cout=0 sum=00110011
* bcd_in1=00000110 bcd_in2=00101000 cout=0 sum=00110100
* bcd_in1=00000110 bcd_in2=00101001 cout=0 sum=00110101
* bcd_in1=00000110 bcd_in2=00110000 cout=0 sum=00110110
* bcd_in1=00000110 bcd_in2=00110001 cout=0 sum=00110111
* bcd_in1=00000110 bcd_in2=00110010 cout=0 sum=00111000
* bcd_in1=00000110 bcd_in2=00110011 cout=0 sum=00111001
* bcd_in1=00000110 bcd_in2=00110100 cout=0 sum=01000000
* bcd_in1=00000110 bcd_in2=00110101 cout=0 sum=01000001
* bcd_in1=00000110 bcd_in2=00110110 cout=0 sum=01000010
* bcd_in1=00000110 bcd_in2=00110111 cout=0 sum=01000011
* bcd_in1=00000110 bcd_in2=00111000 cout=0 sum=01000100
* bcd_in1=00000110 bcd_in2=00111001 cout=0 sum=01000101
* bcd_in1=00000110 bcd_in2=01000000 cout=0 sum=01000110
* bcd_in1=00000110 bcd_in2=01000001 cout=0 sum=01000111
* bcd_in1=00000110 bcd_in2=01000010 cout=0 sum=01001000
* bcd_in1=00000110 bcd_in2=01000011 cout=0 sum=01001001
* bcd_in1=00000110 bcd_in2=01000100 cout=0 sum=01010000
* bcd_in1=00000110 bcd_in2=01000101 cout=0 sum=01010001
* bcd_in1=00000110 bcd_in2=01000110 cout=0 sum=01010010
* bcd_in1=00000110 bcd_in2=01000111 cout=0 sum=01010011
* bcd_in1=00000110 bcd_in2=01001000 cout=0 sum=01010100
* bcd_in1=00000110 bcd_in2=01001001 cout=0 sum=01010101
* bcd_in1=00000110 bcd_in2=01010000 cout=0 sum=01010110
* bcd_in1=00000110 bcd_in2=01010001 cout=0 sum=01010111
* bcd_in1=00000110 bcd_in2=01010010 cout=0 sum=01011000
* bcd_in1=00000110 bcd_in2=01010011 cout=0 sum=01011001
* bcd_in1=00000110 bcd_in2=01010100 cout=0 sum=01100000
* bcd_in1=00000110 bcd_in2=01010101 cout=0 sum=01100001
* bcd_in1=00000110 bcd_in2=01010110 cout=0 sum=01100010
* bcd_in1=00000110 bcd_in2=01010111 cout=0 sum=01100011
* bcd_in1=00000110 bcd_in2=01011000 cout=0 sum=01100100
* bcd_in1=00000110 bcd_in2=01011001 cout=0 sum=01100101
* bcd_in1=00000110 bcd_in2=01100000 cout=0 sum=01100110
* bcd_in1=00000110 bcd_in2=01100001 cout=0 sum=01100111
* bcd_in1=00000110 bcd_in2=01100010 cout=0 sum=01101000
* bcd_in1=00000110 bcd_in2=01100011 cout=0 sum=01101001
* bcd_in1=00000110 bcd_in2=01100100 cout=0 sum=01110000
* bcd_in1=00000110 bcd_in2=01100101 cout=0 sum=01110001
* bcd_in1=00000110 bcd_in2=01100110 cout=0 sum=01110010
* bcd_in1=00000110 bcd_in2=01100111 cout=0 sum=01110011
* bcd_in1=00000110 bcd_in2=01101000 cout=0 sum=01110100
* bcd_in1=00000110 bcd_in2=01101001 cout=0 sum=01110101
* bcd_in1=00000110 bcd_in2=01110000 cout=0 sum=01110110
* bcd_in1=00000110 bcd_in2=01110001 cout=0 sum=01110111
* bcd_in1=00000110 bcd_in2=01110010 cout=0 sum=01111000
* bcd_in1=00000110 bcd_in2=01110011 cout=0 sum=01111001
* bcd_in1=00000110 bcd_in2=01110100 cout=0 sum=10000000
* bcd_in1=00000110 bcd_in2=01110101 cout=0 sum=10000001
* bcd_in1=00000110 bcd_in2=01110110 cout=0 sum=10000010
* bcd_in1=00000110 bcd_in2=01110111 cout=0 sum=10000011
* bcd_in1=00000110 bcd_in2=01111000 cout=0 sum=10000100
* bcd_in1=00000110 bcd_in2=01111001 cout=0 sum=10000101
* bcd_in1=00000110 bcd_in2=10000000 cout=0 sum=10000110
* bcd_in1=00000110 bcd_in2=10000001 cout=0 sum=10000111
* bcd_in1=00000110 bcd_in2=10000010 cout=0 sum=10001000
* bcd_in1=00000110 bcd_in2=10000011 cout=0 sum=10001001
* bcd_in1=00000110 bcd_in2=10000100 cout=0 sum=10010000
* bcd_in1=00000110 bcd_in2=10000101 cout=0 sum=10010001
* bcd_in1=00000110 bcd_in2=10000110 cout=0 sum=10010010
* bcd_in1=00000110 bcd_in2=10000111 cout=0 sum=10010011
* bcd_in1=00000110 bcd_in2=10001000 cout=0 sum=10010100
* bcd_in1=00000110 bcd_in2=10001001 cout=0 sum=10010101
* bcd_in1=00000110 bcd_in2=10010000 cout=0 sum=10010110
* bcd_in1=00000110 bcd_in2=10010001 cout=0 sum=10010111
* bcd_in1=00000110 bcd_in2=10010010 cout=0 sum=10011000
* bcd_in1=00000110 bcd_in2=10010011 cout=0 sum=10011001
* bcd_in1=00000110 bcd_in2=10010100 cout=1 sum=00000000
* bcd_in1=00000110 bcd_in2=10010101 cout=1 sum=00000001
* bcd_in1=00000110 bcd_in2=10010110 cout=1 sum=00000010
* bcd_in1=00000110 bcd_in2=10010111 cout=1 sum=00000011
* bcd_in1=00000110 bcd_in2=10011000 cout=1 sum=00000100
* bcd_in1=00000110 bcd_in2=10011001 cout=1 sum=00000101
* bcd_in1=00000111 bcd_in2=00000000 cout=0 sum=00000111
* bcd_in1=00000111 bcd_in2=00000001 cout=0 sum=00001000
* bcd_in1=00000111 bcd_in2=00000010 cout=0 sum=00001001
* bcd_in1=00000111 bcd_in2=00000011 cout=0 sum=00010000
* bcd_in1=00000111 bcd_in2=00000100 cout=0 sum=00010001
* bcd_in1=00000111 bcd_in2=00000101 cout=0 sum=00010010
* bcd_in1=00000111 bcd_in2=00000110 cout=0 sum=00010011
* bcd_in1=00000111 bcd_in2=00000111 cout=0 sum=00010100
* bcd_in1=00000111 bcd_in2=00001000 cout=0 sum=00010101
* bcd_in1=00000111 bcd_in2=00001001 cout=0 sum=00010110
* bcd_in1=00000111 bcd_in2=00010000 cout=0 sum=00010111
* bcd_in1=00000111 bcd_in2=00010001 cout=0 sum=00011000
* bcd_in1=00000111 bcd_in2=00010010 cout=0 sum=00011001
* bcd_in1=00000111 bcd_in2=00010011 cout=0 sum=00100000
* bcd_in1=00000111 bcd_in2=00010100 cout=0 sum=00100001
* bcd_in1=00000111 bcd_in2=00010101 cout=0 sum=00100010
* bcd_in1=00000111 bcd_in2=00010110 cout=0 sum=00100011
* bcd_in1=00000111 bcd_in2=00010111 cout=0 sum=00100100
* bcd_in1=00000111 bcd_in2=00011000 cout=0 sum=00100101
* bcd_in1=00000111 bcd_in2=00011001 cout=0 sum=00100110
* bcd_in1=00000111 bcd_in2=00100000 cout=0 sum=00100111
* bcd_in1=00000111 bcd_in2=00100001 cout=0 sum=00101000
* bcd_in1=00000111 bcd_in2=00100010 cout=0 sum=00101001
* bcd_in1=00000111 bcd_in2=00100011 cout=0 sum=00110000
* bcd_in1=00000111 bcd_in2=00100100 cout=0 sum=00110001
* bcd_in1=00000111 bcd_in2=00100101 cout=0 sum=00110010
* bcd_in1=00000111 bcd_in2=00100110 cout=0 sum=00110011
* bcd_in1=00000111 bcd_in2=00100111 cout=0 sum=00110100
* bcd_in1=00000111 bcd_in2=00101000 cout=0 sum=00110101
* bcd_in1=00000111 bcd_in2=00101001 cout=0 sum=00110110
* bcd_in1=00000111 bcd_in2=00110000 cout=0 sum=00110111
* bcd_in1=00000111 bcd_in2=00110001 cout=0 sum=00111000
* bcd_in1=00000111 bcd_in2=00110010 cout=0 sum=00111001
* bcd_in1=00000111 bcd_in2=00110011 cout=0 sum=01000000
* bcd_in1=00000111 bcd_in2=00110100 cout=0 sum=01000001
* bcd_in1=00000111 bcd_in2=00110101 cout=0 sum=01000010
* bcd_in1=00000111 bcd_in2=00110110 cout=0 sum=01000011
* bcd_in1=00000111 bcd_in2=00110111 cout=0 sum=01000100
* bcd_in1=00000111 bcd_in2=00111000 cout=0 sum=01000101
* bcd_in1=00000111 bcd_in2=00111001 cout=0 sum=01000110
* bcd_in1=00000111 bcd_in2=01000000 cout=0 sum=01000111
* bcd_in1=00000111 bcd_in2=01000001 cout=0 sum=01001000
* bcd_in1=00000111 bcd_in2=01000010 cout=0 sum=01001001
* bcd_in1=00000111 bcd_in2=01000011 cout=0 sum=01010000
* bcd_in1=00000111 bcd_in2=01000100 cout=0 sum=01010001
* bcd_in1=00000111 bcd_in2=01000101 cout=0 sum=01010010
* bcd_in1=00000111 bcd_in2=01000110 cout=0 sum=01010011
* bcd_in1=00000111 bcd_in2=01000111 cout=0 sum=01010100
* bcd_in1=00000111 bcd_in2=01001000 cout=0 sum=01010101
* bcd_in1=00000111 bcd_in2=01001001 cout=0 sum=01010110
* bcd_in1=00000111 bcd_in2=01010000 cout=0 sum=01010111
* bcd_in1=00000111 bcd_in2=01010001 cout=0 sum=01011000
* bcd_in1=00000111 bcd_in2=01010010 cout=0 sum=01011001
* bcd_in1=00000111 bcd_in2=01010011 cout=0 sum=01100000
* bcd_in1=00000111 bcd_in2=01010100 cout=0 sum=01100001
* bcd_in1=00000111 bcd_in2=01010101 cout=0 sum=01100010
* bcd_in1=00000111 bcd_in2=01010110 cout=0 sum=01100011
* bcd_in1=00000111 bcd_in2=01010111 cout=0 sum=01100100
* bcd_in1=00000111 bcd_in2=01011000 cout=0 sum=01100101
* bcd_in1=00000111 bcd_in2=01011001 cout=0 sum=01100110
* bcd_in1=00000111 bcd_in2=01100000 cout=0 sum=01100111
* bcd_in1=00000111 bcd_in2=01100001 cout=0 sum=01101000
* bcd_in1=00000111 bcd_in2=01100010 cout=0 sum=01101001
* bcd_in1=00000111 bcd_in2=01100011 cout=0 sum=01110000
* bcd_in1=00000111 bcd_in2=01100100 cout=0 sum=01110001
* bcd_in1=00000111 bcd_in2=01100101 cout=0 sum=01110010
* bcd_in1=00000111 bcd_in2=01100110 cout=0 sum=01110011
* bcd_in1=00000111 bcd_in2=01100111 cout=0 sum=01110100
* bcd_in1=00000111 bcd_in2=01101000 cout=0 sum=01110101
* bcd_in1=00000111 bcd_in2=01101001 cout=0 sum=01110110
* bcd_in1=00000111 bcd_in2=01110000 cout=0 sum=01110111
* bcd_in1=00000111 bcd_in2=01110001 cout=0 sum=01111000
* bcd_in1=00000111 bcd_in2=01110010 cout=0 sum=01111001
* bcd_in1=00000111 bcd_in2=01110011 cout=0 sum=10000000
* bcd_in1=00000111 bcd_in2=01110100 cout=0 sum=10000001
* bcd_in1=00000111 bcd_in2=01110101 cout=0 sum=10000010
* bcd_in1=00000111 bcd_in2=01110110 cout=0 sum=10000011
* bcd_in1=00000111 bcd_in2=01110111 cout=0 sum=10000100
* bcd_in1=00000111 bcd_in2=01111000 cout=0 sum=10000101
* bcd_in1=00000111 bcd_in2=01111001 cout=0 sum=10000110
* bcd_in1=00000111 bcd_in2=10000000 cout=0 sum=10000111
* bcd_in1=00000111 bcd_in2=10000001 cout=0 sum=10001000
* bcd_in1=00000111 bcd_in2=10000010 cout=0 sum=10001001
* bcd_in1=00000111 bcd_in2=10000011 cout=0 sum=10010000
* bcd_in1=00000111 bcd_in2=10000100 cout=0 sum=10010001
* bcd_in1=00000111 bcd_in2=10000101 cout=0 sum=10010010
* bcd_in1=00000111 bcd_in2=10000110 cout=0 sum=10010011
* bcd_in1=00000111 bcd_in2=10000111 cout=0 sum=10010100
* bcd_in1=00000111 bcd_in2=10001000 cout=0 sum=10010101
* bcd_in1=00000111 bcd_in2=10001001 cout=0 sum=10010110
* bcd_in1=00000111 bcd_in2=10010000 cout=0 sum=10010111
* bcd_in1=00000111 bcd_in2=10010001 cout=0 sum=10011000
* bcd_in1=00000111 bcd_in2=10010010 cout=0 sum=10011001
* bcd_in1=00000111 bcd_in2=10010011 cout=1 sum=00000000
* bcd_in1=00000111 bcd_in2=10010100 cout=1 sum=00000001
* bcd_in1=00000111 bcd_in2=10010101 cout=1 sum=00000010
* bcd_in1=00000111 bcd_in2=10010110 cout=1 sum=00000011
* bcd_in1=00000111 bcd_in2=10010111 cout=1 sum=00000100
* bcd_in1=00000111 bcd_in2=10011000 cout=1 sum=00000101
* bcd_in1=00000111 bcd_in2=10011001 cout=1 sum=00000110
* bcd_in1=00001000 bcd_in2=00000000 cout=0 sum=00001000
* bcd_in1=00001000 bcd_in2=00000001 cout=0 sum=00001001
* bcd_in1=00001000 bcd_in2=00000010 cout=0 sum=00010000
* bcd_in1=00001000 bcd_in2=00000011 cout=0 sum=00010001
* bcd_in1=00001000 bcd_in2=00000100 cout=0 sum=00010010
* bcd_in1=00001000 bcd_in2=00000101 cout=0 sum=00010011
* bcd_in1=00001000 bcd_in2=00000110 cout=0 sum=00010100
* bcd_in1=00001000 bcd_in2=00000111 cout=0 sum=00010101
* bcd_in1=00001000 bcd_in2=00001000 cout=0 sum=00010110
* bcd_in1=00001000 bcd_in2=00001001 cout=0 sum=00010111
* bcd_in1=00001000 bcd_in2=00010000 cout=0 sum=00011000
* bcd_in1=00001000 bcd_in2=00010001 cout=0 sum=00011001
* bcd_in1=00001000 bcd_in2=00010010 cout=0 sum=00100000
* bcd_in1=00001000 bcd_in2=00010011 cout=0 sum=00100001
* bcd_in1=00001000 bcd_in2=00010100 cout=0 sum=00100010
* bcd_in1=00001000 bcd_in2=00010101 cout=0 sum=00100011
* bcd_in1=00001000 bcd_in2=00010110 cout=0 sum=00100100
* bcd_in1=00001000 bcd_in2=00010111 cout=0 sum=00100101
* bcd_in1=00001000 bcd_in2=00011000 cout=0 sum=00100110
* bcd_in1=00001000 bcd_in2=00011001 cout=0 sum=00100111
* bcd_in1=00001000 bcd_in2=00100000 cout=0 sum=00101000
* bcd_in1=00001000 bcd_in2=00100001 cout=0 sum=00101001
* bcd_in1=00001000 bcd_in2=00100010 cout=0 sum=00110000
* bcd_in1=00001000 bcd_in2=00100011 cout=0 sum=00110001
* bcd_in1=00001000 bcd_in2=00100100 cout=0 sum=00110010
* bcd_in1=00001000 bcd_in2=00100101 cout=0 sum=00110011
* bcd_in1=00001000 bcd_in2=00100110 cout=0 sum=00110100
* bcd_in1=00001000 bcd_in2=00100111 cout=0 sum=00110101
* bcd_in1=00001000 bcd_in2=00101000 cout=0 sum=00110110
* bcd_in1=00001000 bcd_in2=00101001 cout=0 sum=00110111
* bcd_in1=00001000 bcd_in2=00110000 cout=0 sum=00111000
* bcd_in1=00001000 bcd_in2=00110001 cout=0 sum=00111001
* bcd_in1=00001000 bcd_in2=00110010 cout=0 sum=01000000
* bcd_in1=00001000 bcd_in2=00110011 cout=0 sum=01000001
* bcd_in1=00001000 bcd_in2=00110100 cout=0 sum=01000010
* bcd_in1=00001000 bcd_in2=00110101 cout=0 sum=01000011
* bcd_in1=00001000 bcd_in2=00110110 cout=0 sum=01000100
* bcd_in1=00001000 bcd_in2=00110111 cout=0 sum=01000101
* bcd_in1=00001000 bcd_in2=00111000 cout=0 sum=01000110
* bcd_in1=00001000 bcd_in2=00111001 cout=0 sum=01000111
* bcd_in1=00001000 bcd_in2=01000000 cout=0 sum=01001000
* bcd_in1=00001000 bcd_in2=01000001 cout=0 sum=01001001
* bcd_in1=00001000 bcd_in2=01000010 cout=0 sum=01010000
* bcd_in1=00001000 bcd_in2=01000011 cout=0 sum=01010001
* bcd_in1=00001000 bcd_in2=01000100 cout=0 sum=01010010
* bcd_in1=00001000 bcd_in2=01000101 cout=0 sum=01010011
* bcd_in1=00001000 bcd_in2=01000110 cout=0 sum=01010100
* bcd_in1=00001000 bcd_in2=01000111 cout=0 sum=01010101
* bcd_in1=00001000 bcd_in2=01001000 cout=0 sum=01010110
* bcd_in1=00001000 bcd_in2=01001001 cout=0 sum=01010111
* bcd_in1=00001000 bcd_in2=01010000 cout=0 sum=01011000
* bcd_in1=00001000 bcd_in2=01010001 cout=0 sum=01011001
* bcd_in1=00001000 bcd_in2=01010010 cout=0 sum=01100000
* bcd_in1=00001000 bcd_in2=01010011 cout=0 sum=01100001
* bcd_in1=00001000 bcd_in2=01010100 cout=0 sum=01100010
* bcd_in1=00001000 bcd_in2=01010101 cout=0 sum=01100011
* bcd_in1=00001000 bcd_in2=01010110 cout=0 sum=01100100
* bcd_in1=00001000 bcd_in2=01010111 cout=0 sum=01100101
* bcd_in1=00001000 bcd_in2=01011000 cout=0 sum=01100110
* bcd_in1=00001000 bcd_in2=01011001 cout=0 sum=01100111
* bcd_in1=00001000 bcd_in2=01100000 cout=0 sum=01101000
* bcd_in1=00001000 bcd_in2=01100001 cout=0 sum=01101001
* bcd_in1=00001000 bcd_in2=01100010 cout=0 sum=01110000
* bcd_in1=00001000 bcd_in2=01100011 cout=0 sum=01110001
* bcd_in1=00001000 bcd_in2=01100100 cout=0 sum=01110010
* bcd_in1=00001000 bcd_in2=01100101 cout=0 sum=01110011
* bcd_in1=00001000 bcd_in2=01100110 cout=0 sum=01110100
* bcd_in1=00001000 bcd_in2=01100111 cout=0 sum=01110101
* bcd_in1=00001000 bcd_in2=01101000 cout=0 sum=01110110
* bcd_in1=00001000 bcd_in2=01101001 cout=0 sum=01110111
* bcd_in1=00001000 bcd_in2=01110000 cout=0 sum=01111000
* bcd_in1=00001000 bcd_in2=01110001 cout=0 sum=01111001
* bcd_in1=00001000 bcd_in2=01110010 cout=0 sum=10000000
* bcd_in1=00001000 bcd_in2=01110011 cout=0 sum=10000001
* bcd_in1=00001000 bcd_in2=01110100 cout=0 sum=10000010
* bcd_in1=00001000 bcd_in2=01110101 cout=0 sum=10000011
* bcd_in1=00001000 bcd_in2=01110110 cout=0 sum=10000100
* bcd_in1=00001000 bcd_in2=01110111 cout=0 sum=10000101
* bcd_in1=00001000 bcd_in2=01111000 cout=0 sum=10000110
* bcd_in1=00001000 bcd_in2=01111001 cout=0 sum=10000111
* bcd_in1=00001000 bcd_in2=10000000 cout=0 sum=10001000
* bcd_in1=00001000 bcd_in2=10000001 cout=0 sum=10001001
* bcd_in1=00001000 bcd_in2=10000010 cout=0 sum=10010000
* bcd_in1=00001000 bcd_in2=10000011 cout=0 sum=10010001
* bcd_in1=00001000 bcd_in2=10000100 cout=0 sum=10010010
* bcd_in1=00001000 bcd_in2=10000101 cout=0 sum=10010011
* bcd_in1=00001000 bcd_in2=10000110 cout=0 sum=10010100
* bcd_in1=00001000 bcd_in2=10000111 cout=0 sum=10010101
* bcd_in1=00001000 bcd_in2=10001000 cout=0 sum=10010110
* bcd_in1=00001000 bcd_in2=10001001 cout=0 sum=10010111
* bcd_in1=00001000 bcd_in2=10010000 cout=0 sum=10011000
* bcd_in1=00001000 bcd_in2=10010001 cout=0 sum=10011001
* bcd_in1=00001000 bcd_in2=10010010 cout=1 sum=00000000
* bcd_in1=00001000 bcd_in2=10010011 cout=1 sum=00000001
* bcd_in1=00001000 bcd_in2=10010100 cout=1 sum=00000010
* bcd_in1=00001000 bcd_in2=10010101 cout=1 sum=00000011
* bcd_in1=00001000 bcd_in2=10010110 cout=1 sum=00000100
* bcd_in1=00001000 bcd_in2=10010111 cout=1 sum=00000101
* bcd_in1=00001000 bcd_in2=10011000 cout=1 sum=00000110
* bcd_in1=00001000 bcd_in2=10011001 cout=1 sum=00000111
* bcd_in1=00001001 bcd_in2=00000000 cout=0 sum=00001001
* bcd_in1=00001001 bcd_in2=00000001 cout=0 sum=00010000
* bcd_in1=00001001 bcd_in2=00000010 cout=0 sum=00010001
* bcd_in1=00001001 bcd_in2=00000011 cout=0 sum=00010010
* bcd_in1=00001001 bcd_in2=00000100 cout=0 sum=00010011
* bcd_in1=00001001 bcd_in2=00000101 cout=0 sum=00010100
* bcd_in1=00001001 bcd_in2=00000110 cout=0 sum=00010101
* bcd_in1=00001001 bcd_in2=00000111 cout=0 sum=00010110
* bcd_in1=00001001 bcd_in2=00001000 cout=0 sum=00010111
* bcd_in1=00001001 bcd_in2=00001001 cout=0 sum=00011000
* bcd_in1=00001001 bcd_in2=00010000 cout=0 sum=00011001
* bcd_in1=00001001 bcd_in2=00010001 cout=0 sum=00100000
* bcd_in1=00001001 bcd_in2=00010010 cout=0 sum=00100001
* bcd_in1=00001001 bcd_in2=00010011 cout=0 sum=00100010
* bcd_in1=00001001 bcd_in2=00010100 cout=0 sum=00100011
* bcd_in1=00001001 bcd_in2=00010101 cout=0 sum=00100100
* bcd_in1=00001001 bcd_in2=00010110 cout=0 sum=00100101
* bcd_in1=00001001 bcd_in2=00010111 cout=0 sum=00100110
* bcd_in1=00001001 bcd_in2=00011000 cout=0 sum=00100111
* bcd_in1=00001001 bcd_in2=00011001 cout=0 sum=00101000
* bcd_in1=00001001 bcd_in2=00100000 cout=0 sum=00101001
* bcd_in1=00001001 bcd_in2=00100001 cout=0 sum=00110000
* bcd_in1=00001001 bcd_in2=00100010 cout=0 sum=00110001
* bcd_in1=00001001 bcd_in2=00100011 cout=0 sum=00110010
* bcd_in1=00001001 bcd_in2=00100100 cout=0 sum=00110011
* bcd_in1=00001001 bcd_in2=00100101 cout=0 sum=00110100
* bcd_in1=00001001 bcd_in2=00100110 cout=0 sum=00110101
* bcd_in1=00001001 bcd_in2=00100111 cout=0 sum=00110110
* bcd_in1=00001001 bcd_in2=00101000 cout=0 sum=00110111
* bcd_in1=00001001 bcd_in2=00101001 cout=0 sum=00111000
* bcd_in1=00001001 bcd_in2=00110000 cout=0 sum=00111001
* bcd_in1=00001001 bcd_in2=00110001 cout=0 sum=01000000
* bcd_in1=00001001 bcd_in2=00110010 cout=0 sum=01000001
* bcd_in1=00001001 bcd_in2=00110011 cout=0 sum=01000010
* bcd_in1=00001001 bcd_in2=00110100 cout=0 sum=01000011
* bcd_in1=00001001 bcd_in2=00110101 cout=0 sum=01000100
* bcd_in1=00001001 bcd_in2=00110110 cout=0 sum=01000101
* bcd_in1=00001001 bcd_in2=00110111 cout=0 sum=01000110
* bcd_in1=00001001 bcd_in2=00111000 cout=0 sum=01000111
* bcd_in1=00001001 bcd_in2=00111001 cout=0 sum=01001000
* bcd_in1=00001001 bcd_in2=01000000 cout=0 sum=01001001
* bcd_in1=00001001 bcd_in2=01000001 cout=0 sum=01010000
* bcd_in1=00001001 bcd_in2=01000010 cout=0 sum=01010001
* bcd_in1=00001001 bcd_in2=01000011 cout=0 sum=01010010
* bcd_in1=00001001 bcd_in2=01000100 cout=0 sum=01010011
* bcd_in1=00001001 bcd_in2=01000101 cout=0 sum=01010100
* bcd_in1=00001001 bcd_in2=01000110 cout=0 sum=01010101
* bcd_in1=00001001 bcd_in2=01000111 cout=0 sum=01010110
* bcd_in1=00001001 bcd_in2=01001000 cout=0 sum=01010111
* bcd_in1=00001001 bcd_in2=01001001 cout=0 sum=01011000
* bcd_in1=00001001 bcd_in2=01010000 cout=0 sum=01011001
* bcd_in1=00001001 bcd_in2=01010001 cout=0 sum=01100000
* bcd_in1=00001001 bcd_in2=01010010 cout=0 sum=01100001
* bcd_in1=00001001 bcd_in2=01010011 cout=0 sum=01100010
* bcd_in1=00001001 bcd_in2=01010100 cout=0 sum=01100011
* bcd_in1=00001001 bcd_in2=01010101 cout=0 sum=01100100
* bcd_in1=00001001 bcd_in2=01010110 cout=0 sum=01100101
* bcd_in1=00001001 bcd_in2=01010111 cout=0 sum=01100110
* bcd_in1=00001001 bcd_in2=01011000 cout=0 sum=01100111
* bcd_in1=00001001 bcd_in2=01011001 cout=0 sum=01101000
* bcd_in1=00001001 bcd_in2=01100000 cout=0 sum=01101001
* bcd_in1=00001001 bcd_in2=01100001 cout=0 sum=01110000
* bcd_in1=00001001 bcd_in2=01100010 cout=0 sum=01110001
* bcd_in1=00001001 bcd_in2=01100011 cout=0 sum=01110010
* bcd_in1=00001001 bcd_in2=01100100 cout=0 sum=01110011
* bcd_in1=00001001 bcd_in2=01100101 cout=0 sum=01110100
* bcd_in1=00001001 bcd_in2=01100110 cout=0 sum=01110101
* bcd_in1=00001001 bcd_in2=01100111 cout=0 sum=01110110
* bcd_in1=00001001 bcd_in2=01101000 cout=0 sum=01110111
* bcd_in1=00001001 bcd_in2=01101001 cout=0 sum=01111000
* bcd_in1=00001001 bcd_in2=01110000 cout=0 sum=01111001
* bcd_in1=00001001 bcd_in2=01110001 cout=0 sum=10000000
* bcd_in1=00001001 bcd_in2=01110010 cout=0 sum=10000001
* bcd_in1=00001001 bcd_in2=01110011 cout=0 sum=10000010
* bcd_in1=00001001 bcd_in2=01110100 cout=0 sum=10000011
* bcd_in1=00001001 bcd_in2=01110101 cout=0 sum=10000100
* bcd_in1=00001001 bcd_in2=01110110 cout=0 sum=10000101
* bcd_in1=00001001 bcd_in2=01110111 cout=0 sum=10000110
* bcd_in1=00001001 bcd_in2=01111000 cout=0 sum=10000111
* bcd_in1=00001001 bcd_in2=01111001 cout=0 sum=10001000
* bcd_in1=00001001 bcd_in2=10000000 cout=0 sum=10001001
* bcd_in1=00001001 bcd_in2=10000001 cout=0 sum=10010000
* bcd_in1=00001001 bcd_in2=10000010 cout=0 sum=10010001
* bcd_in1=00001001 bcd_in2=10000011 cout=0 sum=10010010
* bcd_in1=00001001 bcd_in2=10000100 cout=0 sum=10010011
* bcd_in1=00001001 bcd_in2=10000101 cout=0 sum=10010100
* bcd_in1=00001001 bcd_in2=10000110 cout=0 sum=10010101
* bcd_in1=00001001 bcd_in2=10000111 cout=0 sum=10010110
* bcd_in1=00001001 bcd_in2=10001000 cout=0 sum=10010111
* bcd_in1=00001001 bcd_in2=10001001 cout=0 sum=10011000
* bcd_in1=00001001 bcd_in2=10010000 cout=0 sum=10011001
* bcd_in1=00001001 bcd_in2=10010001 cout=1 sum=00000000
* bcd_in1=00001001 bcd_in2=10010010 cout=1 sum=00000001
* bcd_in1=00001001 bcd_in2=10010011 cout=1 sum=00000010
* bcd_in1=00001001 bcd_in2=10010100 cout=1 sum=00000011
* bcd_in1=00001001 bcd_in2=10010101 cout=1 sum=00000100
* bcd_in1=00001001 bcd_in2=10010110 cout=1 sum=00000101
* bcd_in1=00001001 bcd_in2=10010111 cout=1 sum=00000110
* bcd_in1=00001001 bcd_in2=10011000 cout=1 sum=00000111
* bcd_in1=00001001 bcd_in2=10011001 cout=1 sum=00001000
* bcd_in1=00010000 bcd_in2=00000000 cout=0 sum=00010000
* bcd_in1=00010000 bcd_in2=00000001 cout=0 sum=00010001
* bcd_in1=00010000 bcd_in2=00000010 cout=0 sum=00010010
* bcd_in1=00010000 bcd_in2=00000011 cout=0 sum=00010011
* bcd_in1=00010000 bcd_in2=00000100 cout=0 sum=00010100
* bcd_in1=00010000 bcd_in2=00000101 cout=0 sum=00010101
* bcd_in1=00010000 bcd_in2=00000110 cout=0 sum=00010110
* bcd_in1=00010000 bcd_in2=00000111 cout=0 sum=00010111
* bcd_in1=00010000 bcd_in2=00001000 cout=0 sum=00011000
* bcd_in1=00010000 bcd_in2=00001001 cout=0 sum=00011001
* bcd_in1=00010000 bcd_in2=00010000 cout=0 sum=00100000
* bcd_in1=00010000 bcd_in2=00010001 cout=0 sum=00100001
* bcd_in1=00010000 bcd_in2=00010010 cout=0 sum=00100010
* bcd_in1=00010000 bcd_in2=00010011 cout=0 sum=00100011
* bcd_in1=00010000 bcd_in2=00010100 cout=0 sum=00100100
* bcd_in1=00010000 bcd_in2=00010101 cout=0 sum=00100101
* bcd_in1=00010000 bcd_in2=00010110 cout=0 sum=00100110
* bcd_in1=00010000 bcd_in2=00010111 cout=0 sum=00100111
* bcd_in1=00010000 bcd_in2=00011000 cout=0 sum=00101000
* bcd_in1=00010000 bcd_in2=00011001 cout=0 sum=00101001
* bcd_in1=00010000 bcd_in2=00100000 cout=0 sum=00110000
* bcd_in1=00010000 bcd_in2=00100001 cout=0 sum=00110001
* bcd_in1=00010000 bcd_in2=00100010 cout=0 sum=00110010
* bcd_in1=00010000 bcd_in2=00100011 cout=0 sum=00110011
* bcd_in1=00010000 bcd_in2=00100100 cout=0 sum=00110100
* bcd_in1=00010000 bcd_in2=00100101 cout=0 sum=00110101
* bcd_in1=00010000 bcd_in2=00100110 cout=0 sum=00110110
* bcd_in1=00010000 bcd_in2=00100111 cout=0 sum=00110111
* bcd_in1=00010000 bcd_in2=00101000 cout=0 sum=00111000
* bcd_in1=00010000 bcd_in2=00101001 cout=0 sum=00111001
* bcd_in1=00010000 bcd_in2=00110000 cout=0 sum=01000000
* bcd_in1=00010000 bcd_in2=00110001 cout=0 sum=01000001
* bcd_in1=00010000 bcd_in2=00110010 cout=0 sum=01000010
* bcd_in1=00010000 bcd_in2=00110011 cout=0 sum=01000011
* bcd_in1=00010000 bcd_in2=00110100 cout=0 sum=01000100
* bcd_in1=00010000 bcd_in2=00110101 cout=0 sum=01000101
* bcd_in1=00010000 bcd_in2=00110110 cout=0 sum=01000110
* bcd_in1=00010000 bcd_in2=00110111 cout=0 sum=01000111
* bcd_in1=00010000 bcd_in2=00111000 cout=0 sum=01001000
* bcd_in1=00010000 bcd_in2=00111001 cout=0 sum=01001001
* bcd_in1=00010000 bcd_in2=01000000 cout=0 sum=01010000
* bcd_in1=00010000 bcd_in2=01000001 cout=0 sum=01010001
* bcd_in1=00010000 bcd_in2=01000010 cout=0 sum=01010010
* bcd_in1=00010000 bcd_in2=01000011 cout=0 sum=01010011
* bcd_in1=00010000 bcd_in2=01000100 cout=0 sum=01010100
* bcd_in1=00010000 bcd_in2=01000101 cout=0 sum=01010101
* bcd_in1=00010000 bcd_in2=01000110 cout=0 sum=01010110
* bcd_in1=00010000 bcd_in2=01000111 cout=0 sum=01010111
* bcd_in1=00010000 bcd_in2=01001000 cout=0 sum=01011000
* bcd_in1=00010000 bcd_in2=01001001 cout=0 sum=01011001
* bcd_in1=00010000 bcd_in2=01010000 cout=0 sum=01100000
* bcd_in1=00010000 bcd_in2=01010001 cout=0 sum=01100001
* bcd_in1=00010000 bcd_in2=01010010 cout=0 sum=01100010
* bcd_in1=00010000 bcd_in2=01010011 cout=0 sum=01100011
* bcd_in1=00010000 bcd_in2=01010100 cout=0 sum=01100100
* bcd_in1=00010000 bcd_in2=01010101 cout=0 sum=01100101
* bcd_in1=00010000 bcd_in2=01010110 cout=0 sum=01100110
* bcd_in1=00010000 bcd_in2=01010111 cout=0 sum=01100111
* bcd_in1=00010000 bcd_in2=01011000 cout=0 sum=01101000
* bcd_in1=00010000 bcd_in2=01011001 cout=0 sum=01101001
* bcd_in1=00010000 bcd_in2=01100000 cout=0 sum=01110000
* bcd_in1=00010000 bcd_in2=01100001 cout=0 sum=01110001
* bcd_in1=00010000 bcd_in2=01100010 cout=0 sum=01110010
* bcd_in1=00010000 bcd_in2=01100011 cout=0 sum=01110011
* bcd_in1=00010000 bcd_in2=01100100 cout=0 sum=01110100
* bcd_in1=00010000 bcd_in2=01100101 cout=0 sum=01110101
* bcd_in1=00010000 bcd_in2=01100110 cout=0 sum=01110110
* bcd_in1=00010000 bcd_in2=01100111 cout=0 sum=01110111
* bcd_in1=00010000 bcd_in2=01101000 cout=0 sum=01111000
* bcd_in1=00010000 bcd_in2=01101001 cout=0 sum=01111001
* bcd_in1=00010000 bcd_in2=01110000 cout=0 sum=10000000
* bcd_in1=00010000 bcd_in2=01110001 cout=0 sum=10000001
* bcd_in1=00010000 bcd_in2=01110010 cout=0 sum=10000010
* bcd_in1=00010000 bcd_in2=01110011 cout=0 sum=10000011
* bcd_in1=00010000 bcd_in2=01110100 cout=0 sum=10000100
* bcd_in1=00010000 bcd_in2=01110101 cout=0 sum=10000101
* bcd_in1=00010000 bcd_in2=01110110 cout=0 sum=10000110
* bcd_in1=00010000 bcd_in2=01110111 cout=0 sum=10000111
* bcd_in1=00010000 bcd_in2=01111000 cout=0 sum=10001000
* bcd_in1=00010000 bcd_in2=01111001 cout=0 sum=10001001
* bcd_in1=00010000 bcd_in2=10000000 cout=0 sum=10010000
* bcd_in1=00010000 bcd_in2=10000001 cout=0 sum=10010001
* bcd_in1=00010000 bcd_in2=10000010 cout=0 sum=10010010
* bcd_in1=00010000 bcd_in2=10000011 cout=0 sum=10010011
* bcd_in1=00010000 bcd_in2=10000100 cout=0 sum=10010100
* bcd_in1=00010000 bcd_in2=10000101 cout=0 sum=10010101
* bcd_in1=00010000 bcd_in2=10000110 cout=0 sum=10010110
* bcd_in1=00010000 bcd_in2=10000111 cout=0 sum=10010111
* bcd_in1=00010000 bcd_in2=10001000 cout=0 sum=10011000
* bcd_in1=00010000 bcd_in2=10001001 cout=0 sum=10011001
* bcd_in1=00010000 bcd_in2=10010000 cout=1 sum=00000000
* bcd_in1=00010000 bcd_in2=10010001 cout=1 sum=00000001
* bcd_in1=00010000 bcd_in2=10010010 cout=1 sum=00000010
* bcd_in1=00010000 bcd_in2=10010011 cout=1 sum=00000011
* bcd_in1=00010000 bcd_in2=10010100 cout=1 sum=00000100
* bcd_in1=00010000 bcd_in2=10010101 cout=1 sum=00000101
* bcd_in1=00010000 bcd_in2=10010110 cout=1 sum=00000110
* bcd_in1=00010000 bcd_in2=10010111 cout=1 sum=00000111
* bcd_in1=00010000 bcd_in2=10011000 cout=1 sum=00001000
* bcd_in1=00010000 bcd_in2=10011001 cout=1 sum=00001001
* bcd_in1=00010001 bcd_in2=00000000 cout=0 sum=00010001
* bcd_in1=00010001 bcd_in2=00000001 cout=0 sum=00010010
* bcd_in1=00010001 bcd_in2=00000010 cout=0 sum=00010011
* bcd_in1=00010001 bcd_in2=00000011 cout=0 sum=00010100
* bcd_in1=00010001 bcd_in2=00000100 cout=0 sum=00010101
* bcd_in1=00010001 bcd_in2=00000101 cout=0 sum=00010110
* bcd_in1=00010001 bcd_in2=00000110 cout=0 sum=00010111
* bcd_in1=00010001 bcd_in2=00000111 cout=0 sum=00011000
* bcd_in1=00010001 bcd_in2=00001000 cout=0 sum=00011001
* bcd_in1=00010001 bcd_in2=00001001 cout=0 sum=00100000
* bcd_in1=00010001 bcd_in2=00010000 cout=0 sum=00100001
* bcd_in1=00010001 bcd_in2=00010001 cout=0 sum=00100010
* bcd_in1=00010001 bcd_in2=00010010 cout=0 sum=00100011
* bcd_in1=00010001 bcd_in2=00010011 cout=0 sum=00100100
* bcd_in1=00010001 bcd_in2=00010100 cout=0 sum=00100101
* bcd_in1=00010001 bcd_in2=00010101 cout=0 sum=00100110
* bcd_in1=00010001 bcd_in2=00010110 cout=0 sum=00100111
* bcd_in1=00010001 bcd_in2=00010111 cout=0 sum=00101000
* bcd_in1=00010001 bcd_in2=00011000 cout=0 sum=00101001
* bcd_in1=00010001 bcd_in2=00011001 cout=0 sum=00110000
* bcd_in1=00010001 bcd_in2=00100000 cout=0 sum=00110001
* bcd_in1=00010001 bcd_in2=00100001 cout=0 sum=00110010
* bcd_in1=00010001 bcd_in2=00100010 cout=0 sum=00110011
* bcd_in1=00010001 bcd_in2=00100011 cout=0 sum=00110100
* bcd_in1=00010001 bcd_in2=00100100 cout=0 sum=00110101
* bcd_in1=00010001 bcd_in2=00100101 cout=0 sum=00110110
* bcd_in1=00010001 bcd_in2=00100110 cout=0 sum=00110111
* bcd_in1=00010001 bcd_in2=00100111 cout=0 sum=00111000
* bcd_in1=00010001 bcd_in2=00101000 cout=0 sum=00111001
* bcd_in1=00010001 bcd_in2=00101001 cout=0 sum=01000000
* bcd_in1=00010001 bcd_in2=00110000 cout=0 sum=01000001
* bcd_in1=00010001 bcd_in2=00110001 cout=0 sum=01000010
* bcd_in1=00010001 bcd_in2=00110010 cout=0 sum=01000011
* bcd_in1=00010001 bcd_in2=00110011 cout=0 sum=01000100
* bcd_in1=00010001 bcd_in2=00110100 cout=0 sum=01000101
* bcd_in1=00010001 bcd_in2=00110101 cout=0 sum=01000110
* bcd_in1=00010001 bcd_in2=00110110 cout=0 sum=01000111
* bcd_in1=00010001 bcd_in2=00110111 cout=0 sum=01001000
* bcd_in1=00010001 bcd_in2=00111000 cout=0 sum=01001001
* bcd_in1=00010001 bcd_in2=00111001 cout=0 sum=01010000
* bcd_in1=00010001 bcd_in2=01000000 cout=0 sum=01010001
* bcd_in1=00010001 bcd_in2=01000001 cout=0 sum=01010010
* bcd_in1=00010001 bcd_in2=01000010 cout=0 sum=01010011
* bcd_in1=00010001 bcd_in2=01000011 cout=0 sum=01010100
* bcd_in1=00010001 bcd_in2=01000100 cout=0 sum=01010101
* bcd_in1=00010001 bcd_in2=01000101 cout=0 sum=01010110
* bcd_in1=00010001 bcd_in2=01000110 cout=0 sum=01010111
* bcd_in1=00010001 bcd_in2=01000111 cout=0 sum=01011000
* bcd_in1=00010001 bcd_in2=01001000 cout=0 sum=01011001
* bcd_in1=00010001 bcd_in2=01001001 cout=0 sum=01100000
* bcd_in1=00010001 bcd_in2=01010000 cout=0 sum=01100001
* bcd_in1=00010001 bcd_in2=01010001 cout=0 sum=01100010
* bcd_in1=00010001 bcd_in2=01010010 cout=0 sum=01100011
* bcd_in1=00010001 bcd_in2=01010011 cout=0 sum=01100100
* bcd_in1=00010001 bcd_in2=01010100 cout=0 sum=01100101
* bcd_in1=00010001 bcd_in2=01010101 cout=0 sum=01100110
* bcd_in1=00010001 bcd_in2=01010110 cout=0 sum=01100111
* bcd_in1=00010001 bcd_in2=01010111 cout=0 sum=01101000
* bcd_in1=00010001 bcd_in2=01011000 cout=0 sum=01101001
* bcd_in1=00010001 bcd_in2=01011001 cout=0 sum=01110000
* bcd_in1=00010001 bcd_in2=01100000 cout=0 sum=01110001
* bcd_in1=00010001 bcd_in2=01100001 cout=0 sum=01110010
* bcd_in1=00010001 bcd_in2=01100010 cout=0 sum=01110011
* bcd_in1=00010001 bcd_in2=01100011 cout=0 sum=01110100
* bcd_in1=00010001 bcd_in2=01100100 cout=0 sum=01110101
* bcd_in1=00010001 bcd_in2=01100101 cout=0 sum=01110110
* bcd_in1=00010001 bcd_in2=01100110 cout=0 sum=01110111
* bcd_in1=00010001 bcd_in2=01100111 cout=0 sum=01111000
* bcd_in1=00010001 bcd_in2=01101000 cout=0 sum=01111001
* bcd_in1=00010001 bcd_in2=01101001 cout=0 sum=10000000
* bcd_in1=00010001 bcd_in2=01110000 cout=0 sum=10000001
* bcd_in1=00010001 bcd_in2=01110001 cout=0 sum=10000010
* bcd_in1=00010001 bcd_in2=01110010 cout=0 sum=10000011
* bcd_in1=00010001 bcd_in2=01110011 cout=0 sum=10000100
* bcd_in1=00010001 bcd_in2=01110100 cout=0 sum=10000101
* bcd_in1=00010001 bcd_in2=01110101 cout=0 sum=10000110
* bcd_in1=00010001 bcd_in2=01110110 cout=0 sum=10000111
* bcd_in1=00010001 bcd_in2=01110111 cout=0 sum=10001000
* bcd_in1=00010001 bcd_in2=01111000 cout=0 sum=10001001
* bcd_in1=00010001 bcd_in2=01111001 cout=0 sum=10010000
* bcd_in1=00010001 bcd_in2=10000000 cout=0 sum=10010001
* bcd_in1=00010001 bcd_in2=10000001 cout=0 sum=10010010
* bcd_in1=00010001 bcd_in2=10000010 cout=0 sum=10010011
* bcd_in1=00010001 bcd_in2=10000011 cout=0 sum=10010100
* bcd_in1=00010001 bcd_in2=10000100 cout=0 sum=10010101
* bcd_in1=00010001 bcd_in2=10000101 cout=0 sum=10010110
* bcd_in1=00010001 bcd_in2=10000110 cout=0 sum=10010111
* bcd_in1=00010001 bcd_in2=10000111 cout=0 sum=10011000
* bcd_in1=00010001 bcd_in2=10001000 cout=0 sum=10011001
* bcd_in1=00010001 bcd_in2=10001001 cout=1 sum=00000000
* bcd_in1=00010001 bcd_in2=10010000 cout=1 sum=00000001
* bcd_in1=00010001 bcd_in2=10010001 cout=1 sum=00000010
* bcd_in1=00010001 bcd_in2=10010010 cout=1 sum=00000011
* bcd_in1=00010001 bcd_in2=10010011 cout=1 sum=00000100
* bcd_in1=00010001 bcd_in2=10010100 cout=1 sum=00000101
* bcd_in1=00010001 bcd_in2=10010101 cout=1 sum=00000110
* bcd_in1=00010001 bcd_in2=10010110 cout=1 sum=00000111
* bcd_in1=00010001 bcd_in2=10010111 cout=1 sum=00001000
* bcd_in1=00010001 bcd_in2=10011000 cout=1 sum=00001001
* bcd_in1=00010001 bcd_in2=10011001 cout=1 sum=00010000
* bcd_in1=00010010 bcd_in2=00000000 cout=0 sum=00010010
* bcd_in1=00010010 bcd_in2=00000001 cout=0 sum=00010011
* bcd_in1=00010010 bcd_in2=00000010 cout=0 sum=00010100
* bcd_in1=00010010 bcd_in2=00000011 cout=0 sum=00010101
* bcd_in1=00010010 bcd_in2=00000100 cout=0 sum=00010110
* bcd_in1=00010010 bcd_in2=00000101 cout=0 sum=00010111
* bcd_in1=00010010 bcd_in2=00000110 cout=0 sum=00011000
* bcd_in1=00010010 bcd_in2=00000111 cout=0 sum=00011001
* bcd_in1=00010010 bcd_in2=00001000 cout=0 sum=00100000
* bcd_in1=00010010 bcd_in2=00001001 cout=0 sum=00100001
* bcd_in1=00010010 bcd_in2=00010000 cout=0 sum=00100010
* bcd_in1=00010010 bcd_in2=00010001 cout=0 sum=00100011
* bcd_in1=00010010 bcd_in2=00010010 cout=0 sum=00100100
* bcd_in1=00010010 bcd_in2=00010011 cout=0 sum=00100101
* bcd_in1=00010010 bcd_in2=00010100 cout=0 sum=00100110
* bcd_in1=00010010 bcd_in2=00010101 cout=0 sum=00100111
* bcd_in1=00010010 bcd_in2=00010110 cout=0 sum=00101000
* bcd_in1=00010010 bcd_in2=00010111 cout=0 sum=00101001
* bcd_in1=00010010 bcd_in2=00011000 cout=0 sum=00110000
* bcd_in1=00010010 bcd_in2=00011001 cout=0 sum=00110001
* bcd_in1=00010010 bcd_in2=00100000 cout=0 sum=00110010
* bcd_in1=00010010 bcd_in2=00100001 cout=0 sum=00110011
* bcd_in1=00010010 bcd_in2=00100010 cout=0 sum=00110100
* bcd_in1=00010010 bcd_in2=00100011 cout=0 sum=00110101
* bcd_in1=00010010 bcd_in2=00100100 cout=0 sum=00110110
* bcd_in1=00010010 bcd_in2=00100101 cout=0 sum=00110111
* bcd_in1=00010010 bcd_in2=00100110 cout=0 sum=00111000
* bcd_in1=00010010 bcd_in2=00100111 cout=0 sum=00111001
* bcd_in1=00010010 bcd_in2=00101000 cout=0 sum=01000000
* bcd_in1=00010010 bcd_in2=00101001 cout=0 sum=01000001
* bcd_in1=00010010 bcd_in2=00110000 cout=0 sum=01000010
* bcd_in1=00010010 bcd_in2=00110001 cout=0 sum=01000011
* bcd_in1=00010010 bcd_in2=00110010 cout=0 sum=01000100
* bcd_in1=00010010 bcd_in2=00110011 cout=0 sum=01000101
* bcd_in1=00010010 bcd_in2=00110100 cout=0 sum=01000110
* bcd_in1=00010010 bcd_in2=00110101 cout=0 sum=01000111
* bcd_in1=00010010 bcd_in2=00110110 cout=0 sum=01001000
* bcd_in1=00010010 bcd_in2=00110111 cout=0 sum=01001001
* bcd_in1=00010010 bcd_in2=00111000 cout=0 sum=01010000
* bcd_in1=00010010 bcd_in2=00111001 cout=0 sum=01010001
* bcd_in1=00010010 bcd_in2=01000000 cout=0 sum=01010010
* bcd_in1=00010010 bcd_in2=01000001 cout=0 sum=01010011
* bcd_in1=00010010 bcd_in2=01000010 cout=0 sum=01010100
* bcd_in1=00010010 bcd_in2=01000011 cout=0 sum=01010101
* bcd_in1=00010010 bcd_in2=01000100 cout=0 sum=01010110
* bcd_in1=00010010 bcd_in2=01000101 cout=0 sum=01010111
* bcd_in1=00010010 bcd_in2=01000110 cout=0 sum=01011000
* bcd_in1=00010010 bcd_in2=01000111 cout=0 sum=01011001
* bcd_in1=00010010 bcd_in2=01001000 cout=0 sum=01100000
* bcd_in1=00010010 bcd_in2=01001001 cout=0 sum=01100001
* bcd_in1=00010010 bcd_in2=01010000 cout=0 sum=01100010
* bcd_in1=00010010 bcd_in2=01010001 cout=0 sum=01100011
* bcd_in1=00010010 bcd_in2=01010010 cout=0 sum=01100100
* bcd_in1=00010010 bcd_in2=01010011 cout=0 sum=01100101
* bcd_in1=00010010 bcd_in2=01010100 cout=0 sum=01100110
* bcd_in1=00010010 bcd_in2=01010101 cout=0 sum=01100111
* bcd_in1=00010010 bcd_in2=01010110 cout=0 sum=01101000
* bcd_in1=00010010 bcd_in2=01010111 cout=0 sum=01101001
* bcd_in1=00010010 bcd_in2=01011000 cout=0 sum=01110000
* bcd_in1=00010010 bcd_in2=01011001 cout=0 sum=01110001
* bcd_in1=00010010 bcd_in2=01100000 cout=0 sum=01110010
* bcd_in1=00010010 bcd_in2=01100001 cout=0 sum=01110011
* bcd_in1=00010010 bcd_in2=01100010 cout=0 sum=01110100
* bcd_in1=00010010 bcd_in2=01100011 cout=0 sum=01110101
* bcd_in1=00010010 bcd_in2=01100100 cout=0 sum=01110110
* bcd_in1=00010010 bcd_in2=01100101 cout=0 sum=01110111
* bcd_in1=00010010 bcd_in2=01100110 cout=0 sum=01111000
* bcd_in1=00010010 bcd_in2=01100111 cout=0 sum=01111001
* bcd_in1=00010010 bcd_in2=01101000 cout=0 sum=10000000
* bcd_in1=00010010 bcd_in2=01101001 cout=0 sum=10000001
* bcd_in1=00010010 bcd_in2=01110000 cout=0 sum=10000010
* bcd_in1=00010010 bcd_in2=01110001 cout=0 sum=10000011
* bcd_in1=00010010 bcd_in2=01110010 cout=0 sum=10000100
* bcd_in1=00010010 bcd_in2=01110011 cout=0 sum=10000101
* bcd_in1=00010010 bcd_in2=01110100 cout=0 sum=10000110
* bcd_in1=00010010 bcd_in2=01110101 cout=0 sum=10000111
* bcd_in1=00010010 bcd_in2=01110110 cout=0 sum=10001000
* bcd_in1=00010010 bcd_in2=01110111 cout=0 sum=10001001
* bcd_in1=00010010 bcd_in2=01111000 cout=0 sum=10010000
* bcd_in1=00010010 bcd_in2=01111001 cout=0 sum=10010001
* bcd_in1=00010010 bcd_in2=10000000 cout=0 sum=10010010
* bcd_in1=00010010 bcd_in2=10000001 cout=0 sum=10010011
* bcd_in1=00010010 bcd_in2=10000010 cout=0 sum=10010100
* bcd_in1=00010010 bcd_in2=10000011 cout=0 sum=10010101
* bcd_in1=00010010 bcd_in2=10000100 cout=0 sum=10010110
* bcd_in1=00010010 bcd_in2=10000101 cout=0 sum=10010111
* bcd_in1=00010010 bcd_in2=10000110 cout=0 sum=10011000
* bcd_in1=00010010 bcd_in2=10000111 cout=0 sum=10011001
* bcd_in1=00010010 bcd_in2=10001000 cout=1 sum=00000000
* bcd_in1=00010010 bcd_in2=10001001 cout=1 sum=00000001
* bcd_in1=00010010 bcd_in2=10010000 cout=1 sum=00000010
* bcd_in1=00010010 bcd_in2=10010001 cout=1 sum=00000011
* bcd_in1=00010010 bcd_in2=10010010 cout=1 sum=00000100
* bcd_in1=00010010 bcd_in2=10010011 cout=1 sum=00000101
* bcd_in1=00010010 bcd_in2=10010100 cout=1 sum=00000110
* bcd_in1=00010010 bcd_in2=10010101 cout=1 sum=00000111
* bcd_in1=00010010 bcd_in2=10010110 cout=1 sum=00001000
* bcd_in1=00010010 bcd_in2=10010111 cout=1 sum=00001001
* bcd_in1=00010010 bcd_in2=10011000 cout=1 sum=00010000
* bcd_in1=00010010 bcd_in2=10011001 cout=1 sum=00010001
* bcd_in1=00010011 bcd_in2=00000000 cout=0 sum=00010011
* bcd_in1=00010011 bcd_in2=00000001 cout=0 sum=00010100
* bcd_in1=00010011 bcd_in2=00000010 cout=0 sum=00010101
* bcd_in1=00010011 bcd_in2=00000011 cout=0 sum=00010110
* bcd_in1=00010011 bcd_in2=00000100 cout=0 sum=00010111
* bcd_in1=00010011 bcd_in2=00000101 cout=0 sum=00011000
* bcd_in1=00010011 bcd_in2=00000110 cout=0 sum=00011001
* bcd_in1=00010011 bcd_in2=00000111 cout=0 sum=00100000
* bcd_in1=00010011 bcd_in2=00001000 cout=0 sum=00100001
* bcd_in1=00010011 bcd_in2=00001001 cout=0 sum=00100010
* bcd_in1=00010011 bcd_in2=00010000 cout=0 sum=00100011
* bcd_in1=00010011 bcd_in2=00010001 cout=0 sum=00100100
* bcd_in1=00010011 bcd_in2=00010010 cout=0 sum=00100101
* bcd_in1=00010011 bcd_in2=00010011 cout=0 sum=00100110
* bcd_in1=00010011 bcd_in2=00010100 cout=0 sum=00100111
* bcd_in1=00010011 bcd_in2=00010101 cout=0 sum=00101000
* bcd_in1=00010011 bcd_in2=00010110 cout=0 sum=00101001
* bcd_in1=00010011 bcd_in2=00010111 cout=0 sum=00110000
* bcd_in1=00010011 bcd_in2=00011000 cout=0 sum=00110001
* bcd_in1=00010011 bcd_in2=00011001 cout=0 sum=00110010
* bcd_in1=00010011 bcd_in2=00100000 cout=0 sum=00110011
* bcd_in1=00010011 bcd_in2=00100001 cout=0 sum=00110100
* bcd_in1=00010011 bcd_in2=00100010 cout=0 sum=00110101
* bcd_in1=00010011 bcd_in2=00100011 cout=0 sum=00110110
* bcd_in1=00010011 bcd_in2=00100100 cout=0 sum=00110111
* bcd_in1=00010011 bcd_in2=00100101 cout=0 sum=00111000
* bcd_in1=00010011 bcd_in2=00100110 cout=0 sum=00111001
* bcd_in1=00010011 bcd_in2=00100111 cout=0 sum=01000000
* bcd_in1=00010011 bcd_in2=00101000 cout=0 sum=01000001
* bcd_in1=00010011 bcd_in2=00101001 cout=0 sum=01000010
* bcd_in1=00010011 bcd_in2=00110000 cout=0 sum=01000011
* bcd_in1=00010011 bcd_in2=00110001 cout=0 sum=01000100
* bcd_in1=00010011 bcd_in2=00110010 cout=0 sum=01000101
* bcd_in1=00010011 bcd_in2=00110011 cout=0 sum=01000110
* bcd_in1=00010011 bcd_in2=00110100 cout=0 sum=01000111
* bcd_in1=00010011 bcd_in2=00110101 cout=0 sum=01001000
* bcd_in1=00010011 bcd_in2=00110110 cout=0 sum=01001001
* bcd_in1=00010011 bcd_in2=00110111 cout=0 sum=01010000
* bcd_in1=00010011 bcd_in2=00111000 cout=0 sum=01010001
* bcd_in1=00010011 bcd_in2=00111001 cout=0 sum=01010010
* bcd_in1=00010011 bcd_in2=01000000 cout=0 sum=01010011
* bcd_in1=00010011 bcd_in2=01000001 cout=0 sum=01010100
* bcd_in1=00010011 bcd_in2=01000010 cout=0 sum=01010101
* bcd_in1=00010011 bcd_in2=01000011 cout=0 sum=01010110
* bcd_in1=00010011 bcd_in2=01000100 cout=0 sum=01010111
* bcd_in1=00010011 bcd_in2=01000101 cout=0 sum=01011000
* bcd_in1=00010011 bcd_in2=01000110 cout=0 sum=01011001
* bcd_in1=00010011 bcd_in2=01000111 cout=0 sum=01100000
* bcd_in1=00010011 bcd_in2=01001000 cout=0 sum=01100001
* bcd_in1=00010011 bcd_in2=01001001 cout=0 sum=01100010
* bcd_in1=00010011 bcd_in2=01010000 cout=0 sum=01100011
* bcd_in1=00010011 bcd_in2=01010001 cout=0 sum=01100100
* bcd_in1=00010011 bcd_in2=01010010 cout=0 sum=01100101
* bcd_in1=00010011 bcd_in2=01010011 cout=0 sum=01100110
* bcd_in1=00010011 bcd_in2=01010100 cout=0 sum=01100111
* bcd_in1=00010011 bcd_in2=01010101 cout=0 sum=01101000
* bcd_in1=00010011 bcd_in2=01010110 cout=0 sum=01101001
* bcd_in1=00010011 bcd_in2=01010111 cout=0 sum=01110000
* bcd_in1=00010011 bcd_in2=01011000 cout=0 sum=01110001
* bcd_in1=00010011 bcd_in2=01011001 cout=0 sum=01110010
* bcd_in1=00010011 bcd_in2=01100000 cout=0 sum=01110011
* bcd_in1=00010011 bcd_in2=01100001 cout=0 sum=01110100
* bcd_in1=00010011 bcd_in2=01100010 cout=0 sum=01110101
* bcd_in1=00010011 bcd_in2=01100011 cout=0 sum=01110110
* bcd_in1=00010011 bcd_in2=01100100 cout=0 sum=01110111
* bcd_in1=00010011 bcd_in2=01100101 cout=0 sum=01111000
* bcd_in1=00010011 bcd_in2=01100110 cout=0 sum=01111001
* bcd_in1=00010011 bcd_in2=01100111 cout=0 sum=10000000
* bcd_in1=00010011 bcd_in2=01101000 cout=0 sum=10000001
* bcd_in1=00010011 bcd_in2=01101001 cout=0 sum=10000010
* bcd_in1=00010011 bcd_in2=01110000 cout=0 sum=10000011
* bcd_in1=00010011 bcd_in2=01110001 cout=0 sum=10000100
* bcd_in1=00010011 bcd_in2=01110010 cout=0 sum=10000101
* bcd_in1=00010011 bcd_in2=01110011 cout=0 sum=10000110
* bcd_in1=00010011 bcd_in2=01110100 cout=0 sum=10000111
* bcd_in1=00010011 bcd_in2=01110101 cout=0 sum=10001000
* bcd_in1=00010011 bcd_in2=01110110 cout=0 sum=10001001
* bcd_in1=00010011 bcd_in2=01110111 cout=0 sum=10010000
* bcd_in1=00010011 bcd_in2=01111000 cout=0 sum=10010001
* bcd_in1=00010011 bcd_in2=01111001 cout=0 sum=10010010
* bcd_in1=00010011 bcd_in2=10000000 cout=0 sum=10010011
* bcd_in1=00010011 bcd_in2=10000001 cout=0 sum=10010100
* bcd_in1=00010011 bcd_in2=10000010 cout=0 sum=10010101
* bcd_in1=00010011 bcd_in2=10000011 cout=0 sum=10010110
* bcd_in1=00010011 bcd_in2=10000100 cout=0 sum=10010111
* bcd_in1=00010011 bcd_in2=10000101 cout=0 sum=10011000
* bcd_in1=00010011 bcd_in2=10000110 cout=0 sum=10011001
* bcd_in1=00010011 bcd_in2=10000111 cout=1 sum=00000000
* bcd_in1=00010011 bcd_in2=10001000 cout=1 sum=00000001
* bcd_in1=00010011 bcd_in2=10001001 cout=1 sum=00000010
* bcd_in1=00010011 bcd_in2=10010000 cout=1 sum=00000011
* bcd_in1=00010011 bcd_in2=10010001 cout=1 sum=00000100
* bcd_in1=00010011 bcd_in2=10010010 cout=1 sum=00000101
* bcd_in1=00010011 bcd_in2=10010011 cout=1 sum=00000110
* bcd_in1=00010011 bcd_in2=10010100 cout=1 sum=00000111
* bcd_in1=00010011 bcd_in2=10010101 cout=1 sum=00001000
* bcd_in1=00010011 bcd_in2=10010110 cout=1 sum=00001001
* bcd_in1=00010011 bcd_in2=10010111 cout=1 sum=00010000
* bcd_in1=00010011 bcd_in2=10011000 cout=1 sum=00010001
* bcd_in1=00010011 bcd_in2=10011001 cout=1 sum=00010010
* bcd_in1=00010100 bcd_in2=00000000 cout=0 sum=00010100
* bcd_in1=00010100 bcd_in2=00000001 cout=0 sum=00010101
* bcd_in1=00010100 bcd_in2=00000010 cout=0 sum=00010110
* bcd_in1=00010100 bcd_in2=00000011 cout=0 sum=00010111
* bcd_in1=00010100 bcd_in2=00000100 cout=0 sum=00011000
* bcd_in1=00010100 bcd_in2=00000101 cout=0 sum=00011001
* bcd_in1=00010100 bcd_in2=00000110 cout=0 sum=00100000
* bcd_in1=00010100 bcd_in2=00000111 cout=0 sum=00100001
* bcd_in1=00010100 bcd_in2=00001000 cout=0 sum=00100010
* bcd_in1=00010100 bcd_in2=00001001 cout=0 sum=00100011
* bcd_in1=00010100 bcd_in2=00010000 cout=0 sum=00100100
* bcd_in1=00010100 bcd_in2=00010001 cout=0 sum=00100101
* bcd_in1=00010100 bcd_in2=00010010 cout=0 sum=00100110
* bcd_in1=00010100 bcd_in2=00010011 cout=0 sum=00100111
* bcd_in1=00010100 bcd_in2=00010100 cout=0 sum=00101000
* bcd_in1=00010100 bcd_in2=00010101 cout=0 sum=00101001
* bcd_in1=00010100 bcd_in2=00010110 cout=0 sum=00110000
* bcd_in1=00010100 bcd_in2=00010111 cout=0 sum=00110001
* bcd_in1=00010100 bcd_in2=00011000 cout=0 sum=00110010
* bcd_in1=00010100 bcd_in2=00011001 cout=0 sum=00110011
* bcd_in1=00010100 bcd_in2=00100000 cout=0 sum=00110100
* bcd_in1=00010100 bcd_in2=00100001 cout=0 sum=00110101
* bcd_in1=00010100 bcd_in2=00100010 cout=0 sum=00110110
* bcd_in1=00010100 bcd_in2=00100011 cout=0 sum=00110111
* bcd_in1=00010100 bcd_in2=00100100 cout=0 sum=00111000
* bcd_in1=00010100 bcd_in2=00100101 cout=0 sum=00111001
* bcd_in1=00010100 bcd_in2=00100110 cout=0 sum=01000000
* bcd_in1=00010100 bcd_in2=00100111 cout=0 sum=01000001
* bcd_in1=00010100 bcd_in2=00101000 cout=0 sum=01000010
* bcd_in1=00010100 bcd_in2=00101001 cout=0 sum=01000011
* bcd_in1=00010100 bcd_in2=00110000 cout=0 sum=01000100
* bcd_in1=00010100 bcd_in2=00110001 cout=0 sum=01000101
* bcd_in1=00010100 bcd_in2=00110010 cout=0 sum=01000110
* bcd_in1=00010100 bcd_in2=00110011 cout=0 sum=01000111
* bcd_in1=00010100 bcd_in2=00110100 cout=0 sum=01001000
* bcd_in1=00010100 bcd_in2=00110101 cout=0 sum=01001001
* bcd_in1=00010100 bcd_in2=00110110 cout=0 sum=01010000
* bcd_in1=00010100 bcd_in2=00110111 cout=0 sum=01010001
* bcd_in1=00010100 bcd_in2=00111000 cout=0 sum=01010010
* bcd_in1=00010100 bcd_in2=00111001 cout=0 sum=01010011
* bcd_in1=00010100 bcd_in2=01000000 cout=0 sum=01010100
* bcd_in1=00010100 bcd_in2=01000001 cout=0 sum=01010101
* bcd_in1=00010100 bcd_in2=01000010 cout=0 sum=01010110
* bcd_in1=00010100 bcd_in2=01000011 cout=0 sum=01010111
* bcd_in1=00010100 bcd_in2=01000100 cout=0 sum=01011000
* bcd_in1=00010100 bcd_in2=01000101 cout=0 sum=01011001
* bcd_in1=00010100 bcd_in2=01000110 cout=0 sum=01100000
* bcd_in1=00010100 bcd_in2=01000111 cout=0 sum=01100001
* bcd_in1=00010100 bcd_in2=01001000 cout=0 sum=01100010
* bcd_in1=00010100 bcd_in2=01001001 cout=0 sum=01100011
* bcd_in1=00010100 bcd_in2=01010000 cout=0 sum=01100100
* bcd_in1=00010100 bcd_in2=01010001 cout=0 sum=01100101
* bcd_in1=00010100 bcd_in2=01010010 cout=0 sum=01100110
* bcd_in1=00010100 bcd_in2=01010011 cout=0 sum=01100111
* bcd_in1=00010100 bcd_in2=01010100 cout=0 sum=01101000
* bcd_in1=00010100 bcd_in2=01010101 cout=0 sum=01101001
* bcd_in1=00010100 bcd_in2=01010110 cout=0 sum=01110000
* bcd_in1=00010100 bcd_in2=01010111 cout=0 sum=01110001
* bcd_in1=00010100 bcd_in2=01011000 cout=0 sum=01110010
* bcd_in1=00010100 bcd_in2=01011001 cout=0 sum=01110011
* bcd_in1=00010100 bcd_in2=01100000 cout=0 sum=01110100
* bcd_in1=00010100 bcd_in2=01100001 cout=0 sum=01110101
* bcd_in1=00010100 bcd_in2=01100010 cout=0 sum=01110110
* bcd_in1=00010100 bcd_in2=01100011 cout=0 sum=01110111
* bcd_in1=00010100 bcd_in2=01100100 cout=0 sum=01111000
* bcd_in1=00010100 bcd_in2=01100101 cout=0 sum=01111001
* bcd_in1=00010100 bcd_in2=01100110 cout=0 sum=10000000
* bcd_in1=00010100 bcd_in2=01100111 cout=0 sum=10000001
* bcd_in1=00010100 bcd_in2=01101000 cout=0 sum=10000010
* bcd_in1=00010100 bcd_in2=01101001 cout=0 sum=10000011
* bcd_in1=00010100 bcd_in2=01110000 cout=0 sum=10000100
* bcd_in1=00010100 bcd_in2=01110001 cout=0 sum=10000101
* bcd_in1=00010100 bcd_in2=01110010 cout=0 sum=10000110
* bcd_in1=00010100 bcd_in2=01110011 cout=0 sum=10000111
* bcd_in1=00010100 bcd_in2=01110100 cout=0 sum=10001000
* bcd_in1=00010100 bcd_in2=01110101 cout=0 sum=10001001
* bcd_in1=00010100 bcd_in2=01110110 cout=0 sum=10010000
* bcd_in1=00010100 bcd_in2=01110111 cout=0 sum=10010001
* bcd_in1=00010100 bcd_in2=01111000 cout=0 sum=10010010
* bcd_in1=00010100 bcd_in2=01111001 cout=0 sum=10010011
* bcd_in1=00010100 bcd_in2=10000000 cout=0 sum=10010100
* bcd_in1=00010100 bcd_in2=10000001 cout=0 sum=10010101
* bcd_in1=00010100 bcd_in2=10000010 cout=0 sum=10010110
* bcd_in1=00010100 bcd_in2=10000011 cout=0 sum=10010111
* bcd_in1=00010100 bcd_in2=10000100 cout=0 sum=10011000
* bcd_in1=00010100 bcd_in2=10000101 cout=0 sum=10011001
* bcd_in1=00010100 bcd_in2=10000110 cout=1 sum=00000000
* bcd_in1=00010100 bcd_in2=10000111 cout=1 sum=00000001
* bcd_in1=00010100 bcd_in2=10001000 cout=1 sum=00000010
* bcd_in1=00010100 bcd_in2=10001001 cout=1 sum=00000011
* bcd_in1=00010100 bcd_in2=10010000 cout=1 sum=00000100
* bcd_in1=00010100 bcd_in2=10010001 cout=1 sum=00000101
* bcd_in1=00010100 bcd_in2=10010010 cout=1 sum=00000110
* bcd_in1=00010100 bcd_in2=10010011 cout=1 sum=00000111
* bcd_in1=00010100 bcd_in2=10010100 cout=1 sum=00001000
* bcd_in1=00010100 bcd_in2=10010101 cout=1 sum=00001001
* bcd_in1=00010100 bcd_in2=10010110 cout=1 sum=00010000
* bcd_in1=00010100 bcd_in2=10010111 cout=1 sum=00010001
* bcd_in1=00010100 bcd_in2=10011000 cout=1 sum=00010010
* bcd_in1=00010100 bcd_in2=10011001 cout=1 sum=00010011
* bcd_in1=00010101 bcd_in2=00000000 cout=0 sum=00010101
* bcd_in1=00010101 bcd_in2=00000001 cout=0 sum=00010110
* bcd_in1=00010101 bcd_in2=00000010 cout=0 sum=00010111
* bcd_in1=00010101 bcd_in2=00000011 cout=0 sum=00011000
* bcd_in1=00010101 bcd_in2=00000100 cout=0 sum=00011001
* bcd_in1=00010101 bcd_in2=00000101 cout=0 sum=00100000
* bcd_in1=00010101 bcd_in2=00000110 cout=0 sum=00100001
* bcd_in1=00010101 bcd_in2=00000111 cout=0 sum=00100010
* bcd_in1=00010101 bcd_in2=00001000 cout=0 sum=00100011
* bcd_in1=00010101 bcd_in2=00001001 cout=0 sum=00100100
* bcd_in1=00010101 bcd_in2=00010000 cout=0 sum=00100101
* bcd_in1=00010101 bcd_in2=00010001 cout=0 sum=00100110
* bcd_in1=00010101 bcd_in2=00010010 cout=0 sum=00100111
* bcd_in1=00010101 bcd_in2=00010011 cout=0 sum=00101000
* bcd_in1=00010101 bcd_in2=00010100 cout=0 sum=00101001
* bcd_in1=00010101 bcd_in2=00010101 cout=0 sum=00110000
* bcd_in1=00010101 bcd_in2=00010110 cout=0 sum=00110001
* bcd_in1=00010101 bcd_in2=00010111 cout=0 sum=00110010
* bcd_in1=00010101 bcd_in2=00011000 cout=0 sum=00110011
* bcd_in1=00010101 bcd_in2=00011001 cout=0 sum=00110100
* bcd_in1=00010101 bcd_in2=00100000 cout=0 sum=00110101
* bcd_in1=00010101 bcd_in2=00100001 cout=0 sum=00110110
* bcd_in1=00010101 bcd_in2=00100010 cout=0 sum=00110111
* bcd_in1=00010101 bcd_in2=00100011 cout=0 sum=00111000
* bcd_in1=00010101 bcd_in2=00100100 cout=0 sum=00111001
* bcd_in1=00010101 bcd_in2=00100101 cout=0 sum=01000000
* bcd_in1=00010101 bcd_in2=00100110 cout=0 sum=01000001
* bcd_in1=00010101 bcd_in2=00100111 cout=0 sum=01000010
* bcd_in1=00010101 bcd_in2=00101000 cout=0 sum=01000011
* bcd_in1=00010101 bcd_in2=00101001 cout=0 sum=01000100
* bcd_in1=00010101 bcd_in2=00110000 cout=0 sum=01000101
* bcd_in1=00010101 bcd_in2=00110001 cout=0 sum=01000110
* bcd_in1=00010101 bcd_in2=00110010 cout=0 sum=01000111
* bcd_in1=00010101 bcd_in2=00110011 cout=0 sum=01001000
* bcd_in1=00010101 bcd_in2=00110100 cout=0 sum=01001001
* bcd_in1=00010101 bcd_in2=00110101 cout=0 sum=01010000
* bcd_in1=00010101 bcd_in2=00110110 cout=0 sum=01010001
* bcd_in1=00010101 bcd_in2=00110111 cout=0 sum=01010010
* bcd_in1=00010101 bcd_in2=00111000 cout=0 sum=01010011
* bcd_in1=00010101 bcd_in2=00111001 cout=0 sum=01010100
* bcd_in1=00010101 bcd_in2=01000000 cout=0 sum=01010101
* bcd_in1=00010101 bcd_in2=01000001 cout=0 sum=01010110
* bcd_in1=00010101 bcd_in2=01000010 cout=0 sum=01010111
* bcd_in1=00010101 bcd_in2=01000011 cout=0 sum=01011000
* bcd_in1=00010101 bcd_in2=01000100 cout=0 sum=01011001
* bcd_in1=00010101 bcd_in2=01000101 cout=0 sum=01100000
* bcd_in1=00010101 bcd_in2=01000110 cout=0 sum=01100001
* bcd_in1=00010101 bcd_in2=01000111 cout=0 sum=01100010
* bcd_in1=00010101 bcd_in2=01001000 cout=0 sum=01100011
* bcd_in1=00010101 bcd_in2=01001001 cout=0 sum=01100100
* bcd_in1=00010101 bcd_in2=01010000 cout=0 sum=01100101
* bcd_in1=00010101 bcd_in2=01010001 cout=0 sum=01100110
* bcd_in1=00010101 bcd_in2=01010010 cout=0 sum=01100111
* bcd_in1=00010101 bcd_in2=01010011 cout=0 sum=01101000
* bcd_in1=00010101 bcd_in2=01010100 cout=0 sum=01101001
* bcd_in1=00010101 bcd_in2=01010101 cout=0 sum=01110000
* bcd_in1=00010101 bcd_in2=01010110 cout=0 sum=01110001
* bcd_in1=00010101 bcd_in2=01010111 cout=0 sum=01110010
* bcd_in1=00010101 bcd_in2=01011000 cout=0 sum=01110011
* bcd_in1=00010101 bcd_in2=01011001 cout=0 sum=01110100
* bcd_in1=00010101 bcd_in2=01100000 cout=0 sum=01110101
* bcd_in1=00010101 bcd_in2=01100001 cout=0 sum=01110110
* bcd_in1=00010101 bcd_in2=01100010 cout=0 sum=01110111
* bcd_in1=00010101 bcd_in2=01100011 cout=0 sum=01111000
* bcd_in1=00010101 bcd_in2=01100100 cout=0 sum=01111001
* bcd_in1=00010101 bcd_in2=01100101 cout=0 sum=10000000
* bcd_in1=00010101 bcd_in2=01100110 cout=0 sum=10000001
* bcd_in1=00010101 bcd_in2=01100111 cout=0 sum=10000010
* bcd_in1=00010101 bcd_in2=01101000 cout=0 sum=10000011
* bcd_in1=00010101 bcd_in2=01101001 cout=0 sum=10000100
* bcd_in1=00010101 bcd_in2=01110000 cout=0 sum=10000101
* bcd_in1=00010101 bcd_in2=01110001 cout=0 sum=10000110
* bcd_in1=00010101 bcd_in2=01110010 cout=0 sum=10000111
* bcd_in1=00010101 bcd_in2=01110011 cout=0 sum=10001000
* bcd_in1=00010101 bcd_in2=01110100 cout=0 sum=10001001
* bcd_in1=00010101 bcd_in2=01110101 cout=0 sum=10010000
* bcd_in1=00010101 bcd_in2=01110110 cout=0 sum=10010001
* bcd_in1=00010101 bcd_in2=01110111 cout=0 sum=10010010
* bcd_in1=00010101 bcd_in2=01111000 cout=0 sum=10010011
* bcd_in1=00010101 bcd_in2=01111001 cout=0 sum=10010100
* bcd_in1=00010101 bcd_in2=10000000 cout=0 sum=10010101
* bcd_in1=00010101 bcd_in2=10000001 cout=0 sum=10010110
* bcd_in1=00010101 bcd_in2=10000010 cout=0 sum=10010111
* bcd_in1=00010101 bcd_in2=10000011 cout=0 sum=10011000
* bcd_in1=00010101 bcd_in2=10000100 cout=0 sum=10011001
* bcd_in1=00010101 bcd_in2=10000101 cout=1 sum=00000000
* bcd_in1=00010101 bcd_in2=10000110 cout=1 sum=00000001
* bcd_in1=00010101 bcd_in2=10000111 cout=1 sum=00000010
* bcd_in1=00010101 bcd_in2=10001000 cout=1 sum=00000011
* bcd_in1=00010101 bcd_in2=10001001 cout=1 sum=00000100
* bcd_in1=00010101 bcd_in2=10010000 cout=1 sum=00000101
* bcd_in1=00010101 bcd_in2=10010001 cout=1 sum=00000110
* bcd_in1=00010101 bcd_in2=10010010 cout=1 sum=00000111
* bcd_in1=00010101 bcd_in2=10010011 cout=1 sum=00001000
* bcd_in1=00010101 bcd_in2=10010100 cout=1 sum=00001001
* bcd_in1=00010101 bcd_in2=10010101 cout=1 sum=00010000
* bcd_in1=00010101 bcd_in2=10010110 cout=1 sum=00010001
* bcd_in1=00010101 bcd_in2=10010111 cout=1 sum=00010010
* bcd_in1=00010101 bcd_in2=10011000 cout=1 sum=00010011
* bcd_in1=00010101 bcd_in2=10011001 cout=1 sum=00010100
* bcd_in1=00010110 bcd_in2=00000000 cout=0 sum=00010110
* bcd_in1=00010110 bcd_in2=00000001 cout=0 sum=00010111
* bcd_in1=00010110 bcd_in2=00000010 cout=0 sum=00011000
* bcd_in1=00010110 bcd_in2=00000011 cout=0 sum=00011001
* bcd_in1=00010110 bcd_in2=00000100 cout=0 sum=00100000
* bcd_in1=00010110 bcd_in2=00000101 cout=0 sum=00100001
* bcd_in1=00010110 bcd_in2=00000110 cout=0 sum=00100010
* bcd_in1=00010110 bcd_in2=00000111 cout=0 sum=00100011
* bcd_in1=00010110 bcd_in2=00001000 cout=0 sum=00100100
* bcd_in1=00010110 bcd_in2=00001001 cout=0 sum=00100101
* bcd_in1=00010110 bcd_in2=00010000 cout=0 sum=00100110
* bcd_in1=00010110 bcd_in2=00010001 cout=0 sum=00100111
* bcd_in1=00010110 bcd_in2=00010010 cout=0 sum=00101000
* bcd_in1=00010110 bcd_in2=00010011 cout=0 sum=00101001
* bcd_in1=00010110 bcd_in2=00010100 cout=0 sum=00110000
* bcd_in1=00010110 bcd_in2=00010101 cout=0 sum=00110001
* bcd_in1=00010110 bcd_in2=00010110 cout=0 sum=00110010
* bcd_in1=00010110 bcd_in2=00010111 cout=0 sum=00110011
* bcd_in1=00010110 bcd_in2=00011000 cout=0 sum=00110100
* bcd_in1=00010110 bcd_in2=00011001 cout=0 sum=00110101
* bcd_in1=00010110 bcd_in2=00100000 cout=0 sum=00110110
* bcd_in1=00010110 bcd_in2=00100001 cout=0 sum=00110111
* bcd_in1=00010110 bcd_in2=00100010 cout=0 sum=00111000
* bcd_in1=00010110 bcd_in2=00100011 cout=0 sum=00111001
* bcd_in1=00010110 bcd_in2=00100100 cout=0 sum=01000000
* bcd_in1=00010110 bcd_in2=00100101 cout=0 sum=01000001
* bcd_in1=00010110 bcd_in2=00100110 cout=0 sum=01000010
* bcd_in1=00010110 bcd_in2=00100111 cout=0 sum=01000011
* bcd_in1=00010110 bcd_in2=00101000 cout=0 sum=01000100
* bcd_in1=00010110 bcd_in2=00101001 cout=0 sum=01000101
* bcd_in1=00010110 bcd_in2=00110000 cout=0 sum=01000110
* bcd_in1=00010110 bcd_in2=00110001 cout=0 sum=01000111
* bcd_in1=00010110 bcd_in2=00110010 cout=0 sum=01001000
* bcd_in1=00010110 bcd_in2=00110011 cout=0 sum=01001001
* bcd_in1=00010110 bcd_in2=00110100 cout=0 sum=01010000
* bcd_in1=00010110 bcd_in2=00110101 cout=0 sum=01010001
* bcd_in1=00010110 bcd_in2=00110110 cout=0 sum=01010010
* bcd_in1=00010110 bcd_in2=00110111 cout=0 sum=01010011
* bcd_in1=00010110 bcd_in2=00111000 cout=0 sum=01010100
* bcd_in1=00010110 bcd_in2=00111001 cout=0 sum=01010101
* bcd_in1=00010110 bcd_in2=01000000 cout=0 sum=01010110
* bcd_in1=00010110 bcd_in2=01000001 cout=0 sum=01010111
* bcd_in1=00010110 bcd_in2=01000010 cout=0 sum=01011000
* bcd_in1=00010110 bcd_in2=01000011 cout=0 sum=01011001
* bcd_in1=00010110 bcd_in2=01000100 cout=0 sum=01100000
* bcd_in1=00010110 bcd_in2=01000101 cout=0 sum=01100001
* bcd_in1=00010110 bcd_in2=01000110 cout=0 sum=01100010
* bcd_in1=00010110 bcd_in2=01000111 cout=0 sum=01100011
* bcd_in1=00010110 bcd_in2=01001000 cout=0 sum=01100100
* bcd_in1=00010110 bcd_in2=01001001 cout=0 sum=01100101
* bcd_in1=00010110 bcd_in2=01010000 cout=0 sum=01100110
* bcd_in1=00010110 bcd_in2=01010001 cout=0 sum=01100111
* bcd_in1=00010110 bcd_in2=01010010 cout=0 sum=01101000
* bcd_in1=00010110 bcd_in2=01010011 cout=0 sum=01101001
* bcd_in1=00010110 bcd_in2=01010100 cout=0 sum=01110000
* bcd_in1=00010110 bcd_in2=01010101 cout=0 sum=01110001
* bcd_in1=00010110 bcd_in2=01010110 cout=0 sum=01110010
* bcd_in1=00010110 bcd_in2=01010111 cout=0 sum=01110011
* bcd_in1=00010110 bcd_in2=01011000 cout=0 sum=01110100
* bcd_in1=00010110 bcd_in2=01011001 cout=0 sum=01110101
* bcd_in1=00010110 bcd_in2=01100000 cout=0 sum=01110110
* bcd_in1=00010110 bcd_in2=01100001 cout=0 sum=01110111
* bcd_in1=00010110 bcd_in2=01100010 cout=0 sum=01111000
* bcd_in1=00010110 bcd_in2=01100011 cout=0 sum=01111001
* bcd_in1=00010110 bcd_in2=01100100 cout=0 sum=10000000
* bcd_in1=00010110 bcd_in2=01100101 cout=0 sum=10000001
* bcd_in1=00010110 bcd_in2=01100110 cout=0 sum=10000010
* bcd_in1=00010110 bcd_in2=01100111 cout=0 sum=10000011
* bcd_in1=00010110 bcd_in2=01101000 cout=0 sum=10000100
* bcd_in1=00010110 bcd_in2=01101001 cout=0 sum=10000101
* bcd_in1=00010110 bcd_in2=01110000 cout=0 sum=10000110
* bcd_in1=00010110 bcd_in2=01110001 cout=0 sum=10000111
* bcd_in1=00010110 bcd_in2=01110010 cout=0 sum=10001000
* bcd_in1=00010110 bcd_in2=01110011 cout=0 sum=10001001
* bcd_in1=00010110 bcd_in2=01110100 cout=0 sum=10010000
* bcd_in1=00010110 bcd_in2=01110101 cout=0 sum=10010001
* bcd_in1=00010110 bcd_in2=01110110 cout=0 sum=10010010
* bcd_in1=00010110 bcd_in2=01110111 cout=0 sum=10010011
* bcd_in1=00010110 bcd_in2=01111000 cout=0 sum=10010100
* bcd_in1=00010110 bcd_in2=01111001 cout=0 sum=10010101
* bcd_in1=00010110 bcd_in2=10000000 cout=0 sum=10010110
* bcd_in1=00010110 bcd_in2=10000001 cout=0 sum=10010111
* bcd_in1=00010110 bcd_in2=10000010 cout=0 sum=10011000
* bcd_in1=00010110 bcd_in2=10000011 cout=0 sum=10011001
* bcd_in1=00010110 bcd_in2=10000100 cout=1 sum=00000000
* bcd_in1=00010110 bcd_in2=10000101 cout=1 sum=00000001
* bcd_in1=00010110 bcd_in2=10000110 cout=1 sum=00000010
* bcd_in1=00010110 bcd_in2=10000111 cout=1 sum=00000011
* bcd_in1=00010110 bcd_in2=10001000 cout=1 sum=00000100
* bcd_in1=00010110 bcd_in2=10001001 cout=1 sum=00000101
* bcd_in1=00010110 bcd_in2=10010000 cout=1 sum=00000110
* bcd_in1=00010110 bcd_in2=10010001 cout=1 sum=00000111
* bcd_in1=00010110 bcd_in2=10010010 cout=1 sum=00001000
* bcd_in1=00010110 bcd_in2=10010011 cout=1 sum=00001001
* bcd_in1=00010110 bcd_in2=10010100 cout=1 sum=00010000
* bcd_in1=00010110 bcd_in2=10010101 cout=1 sum=00010001
* bcd_in1=00010110 bcd_in2=10010110 cout=1 sum=00010010
* bcd_in1=00010110 bcd_in2=10010111 cout=1 sum=00010011
* bcd_in1=00010110 bcd_in2=10011000 cout=1 sum=00010100
* bcd_in1=00010110 bcd_in2=10011001 cout=1 sum=00010101
* bcd_in1=00010111 bcd_in2=00000000 cout=0 sum=00010111
* bcd_in1=00010111 bcd_in2=00000001 cout=0 sum=00011000
* bcd_in1=00010111 bcd_in2=00000010 cout=0 sum=00011001
* bcd_in1=00010111 bcd_in2=00000011 cout=0 sum=00100000
* bcd_in1=00010111 bcd_in2=00000100 cout=0 sum=00100001
* bcd_in1=00010111 bcd_in2=00000101 cout=0 sum=00100010
* bcd_in1=00010111 bcd_in2=00000110 cout=0 sum=00100011
* bcd_in1=00010111 bcd_in2=00000111 cout=0 sum=00100100
* bcd_in1=00010111 bcd_in2=00001000 cout=0 sum=00100101
* bcd_in1=00010111 bcd_in2=00001001 cout=0 sum=00100110
* bcd_in1=00010111 bcd_in2=00010000 cout=0 sum=00100111
* bcd_in1=00010111 bcd_in2=00010001 cout=0 sum=00101000
* bcd_in1=00010111 bcd_in2=00010010 cout=0 sum=00101001
* bcd_in1=00010111 bcd_in2=00010011 cout=0 sum=00110000
* bcd_in1=00010111 bcd_in2=00010100 cout=0 sum=00110001
* bcd_in1=00010111 bcd_in2=00010101 cout=0 sum=00110010
* bcd_in1=00010111 bcd_in2=00010110 cout=0 sum=00110011
* bcd_in1=00010111 bcd_in2=00010111 cout=0 sum=00110100
* bcd_in1=00010111 bcd_in2=00011000 cout=0 sum=00110101
* bcd_in1=00010111 bcd_in2=00011001 cout=0 sum=00110110
* bcd_in1=00010111 bcd_in2=00100000 cout=0 sum=00110111
* bcd_in1=00010111 bcd_in2=00100001 cout=0 sum=00111000
* bcd_in1=00010111 bcd_in2=00100010 cout=0 sum=00111001
* bcd_in1=00010111 bcd_in2=00100011 cout=0 sum=01000000
* bcd_in1=00010111 bcd_in2=00100100 cout=0 sum=01000001
* bcd_in1=00010111 bcd_in2=00100101 cout=0 sum=01000010
* bcd_in1=00010111 bcd_in2=00100110 cout=0 sum=01000011
* bcd_in1=00010111 bcd_in2=00100111 cout=0 sum=01000100
* bcd_in1=00010111 bcd_in2=00101000 cout=0 sum=01000101
* bcd_in1=00010111 bcd_in2=00101001 cout=0 sum=01000110
* bcd_in1=00010111 bcd_in2=00110000 cout=0 sum=01000111
* bcd_in1=00010111 bcd_in2=00110001 cout=0 sum=01001000
* bcd_in1=00010111 bcd_in2=00110010 cout=0 sum=01001001
* bcd_in1=00010111 bcd_in2=00110011 cout=0 sum=01010000
* bcd_in1=00010111 bcd_in2=00110100 cout=0 sum=01010001
* bcd_in1=00010111 bcd_in2=00110101 cout=0 sum=01010010
* bcd_in1=00010111 bcd_in2=00110110 cout=0 sum=01010011
* bcd_in1=00010111 bcd_in2=00110111 cout=0 sum=01010100
* bcd_in1=00010111 bcd_in2=00111000 cout=0 sum=01010101
* bcd_in1=00010111 bcd_in2=00111001 cout=0 sum=01010110
* bcd_in1=00010111 bcd_in2=01000000 cout=0 sum=01010111
* bcd_in1=00010111 bcd_in2=01000001 cout=0 sum=01011000
* bcd_in1=00010111 bcd_in2=01000010 cout=0 sum=01011001
* bcd_in1=00010111 bcd_in2=01000011 cout=0 sum=01100000
* bcd_in1=00010111 bcd_in2=01000100 cout=0 sum=01100001
* bcd_in1=00010111 bcd_in2=01000101 cout=0 sum=01100010
* bcd_in1=00010111 bcd_in2=01000110 cout=0 sum=01100011
* bcd_in1=00010111 bcd_in2=01000111 cout=0 sum=01100100
* bcd_in1=00010111 bcd_in2=01001000 cout=0 sum=01100101
* bcd_in1=00010111 bcd_in2=01001001 cout=0 sum=01100110
* bcd_in1=00010111 bcd_in2=01010000 cout=0 sum=01100111
* bcd_in1=00010111 bcd_in2=01010001 cout=0 sum=01101000
* bcd_in1=00010111 bcd_in2=01010010 cout=0 sum=01101001
* bcd_in1=00010111 bcd_in2=01010011 cout=0 sum=01110000
* bcd_in1=00010111 bcd_in2=01010100 cout=0 sum=01110001
* bcd_in1=00010111 bcd_in2=01010101 cout=0 sum=01110010
* bcd_in1=00010111 bcd_in2=01010110 cout=0 sum=01110011
* bcd_in1=00010111 bcd_in2=01010111 cout=0 sum=01110100
* bcd_in1=00010111 bcd_in2=01011000 cout=0 sum=01110101
* bcd_in1=00010111 bcd_in2=01011001 cout=0 sum=01110110
* bcd_in1=00010111 bcd_in2=01100000 cout=0 sum=01110111
* bcd_in1=00010111 bcd_in2=01100001 cout=0 sum=01111000
* bcd_in1=00010111 bcd_in2=01100010 cout=0 sum=01111001
* bcd_in1=00010111 bcd_in2=01100011 cout=0 sum=10000000
* bcd_in1=00010111 bcd_in2=01100100 cout=0 sum=10000001
* bcd_in1=00010111 bcd_in2=01100101 cout=0 sum=10000010
* bcd_in1=00010111 bcd_in2=01100110 cout=0 sum=10000011
* bcd_in1=00010111 bcd_in2=01100111 cout=0 sum=10000100
* bcd_in1=00010111 bcd_in2=01101000 cout=0 sum=10000101
* bcd_in1=00010111 bcd_in2=01101001 cout=0 sum=10000110
* bcd_in1=00010111 bcd_in2=01110000 cout=0 sum=10000111
* bcd_in1=00010111 bcd_in2=01110001 cout=0 sum=10001000
* bcd_in1=00010111 bcd_in2=01110010 cout=0 sum=10001001
* bcd_in1=00010111 bcd_in2=01110011 cout=0 sum=10010000
* bcd_in1=00010111 bcd_in2=01110100 cout=0 sum=10010001
* bcd_in1=00010111 bcd_in2=01110101 cout=0 sum=10010010
* bcd_in1=00010111 bcd_in2=01110110 cout=0 sum=10010011
* bcd_in1=00010111 bcd_in2=01110111 cout=0 sum=10010100
* bcd_in1=00010111 bcd_in2=01111000 cout=0 sum=10010101
* bcd_in1=00010111 bcd_in2=01111001 cout=0 sum=10010110
* bcd_in1=00010111 bcd_in2=10000000 cout=0 sum=10010111
* bcd_in1=00010111 bcd_in2=10000001 cout=0 sum=10011000
* bcd_in1=00010111 bcd_in2=10000010 cout=0 sum=10011001
* bcd_in1=00010111 bcd_in2=10000011 cout=1 sum=00000000
* bcd_in1=00010111 bcd_in2=10000100 cout=1 sum=00000001
* bcd_in1=00010111 bcd_in2=10000101 cout=1 sum=00000010
* bcd_in1=00010111 bcd_in2=10000110 cout=1 sum=00000011
* bcd_in1=00010111 bcd_in2=10000111 cout=1 sum=00000100
* bcd_in1=00010111 bcd_in2=10001000 cout=1 sum=00000101
* bcd_in1=00010111 bcd_in2=10001001 cout=1 sum=00000110
* bcd_in1=00010111 bcd_in2=10010000 cout=1 sum=00000111
* bcd_in1=00010111 bcd_in2=10010001 cout=1 sum=00001000
* bcd_in1=00010111 bcd_in2=10010010 cout=1 sum=00001001
* bcd_in1=00010111 bcd_in2=10010011 cout=1 sum=00010000
* bcd_in1=00010111 bcd_in2=10010100 cout=1 sum=00010001
* bcd_in1=00010111 bcd_in2=10010101 cout=1 sum=00010010
* bcd_in1=00010111 bcd_in2=10010110 cout=1 sum=00010011
* bcd_in1=00010111 bcd_in2=10010111 cout=1 sum=00010100
* bcd_in1=00010111 bcd_in2=10011000 cout=1 sum=00010101
* bcd_in1=00010111 bcd_in2=10011001 cout=1 sum=00010110
* bcd_in1=00011000 bcd_in2=00000000 cout=0 sum=00011000
* bcd_in1=00011000 bcd_in2=00000001 cout=0 sum=00011001
* bcd_in1=00011000 bcd_in2=00000010 cout=0 sum=00100000
* bcd_in1=00011000 bcd_in2=00000011 cout=0 sum=00100001
* bcd_in1=00011000 bcd_in2=00000100 cout=0 sum=00100010
* bcd_in1=00011000 bcd_in2=00000101 cout=0 sum=00100011
* bcd_in1=00011000 bcd_in2=00000110 cout=0 sum=00100100
* bcd_in1=00011000 bcd_in2=00000111 cout=0 sum=00100101
* bcd_in1=00011000 bcd_in2=00001000 cout=0 sum=00100110
* bcd_in1=00011000 bcd_in2=00001001 cout=0 sum=00100111
* bcd_in1=00011000 bcd_in2=00010000 cout=0 sum=00101000
* bcd_in1=00011000 bcd_in2=00010001 cout=0 sum=00101001
* bcd_in1=00011000 bcd_in2=00010010 cout=0 sum=00110000
* bcd_in1=00011000 bcd_in2=00010011 cout=0 sum=00110001
* bcd_in1=00011000 bcd_in2=00010100 cout=0 sum=00110010
* bcd_in1=00011000 bcd_in2=00010101 cout=0 sum=00110011
* bcd_in1=00011000 bcd_in2=00010110 cout=0 sum=00110100
* bcd_in1=00011000 bcd_in2=00010111 cout=0 sum=00110101
* bcd_in1=00011000 bcd_in2=00011000 cout=0 sum=00110110
* bcd_in1=00011000 bcd_in2=00011001 cout=0 sum=00110111
* bcd_in1=00011000 bcd_in2=00100000 cout=0 sum=00111000
* bcd_in1=00011000 bcd_in2=00100001 cout=0 sum=00111001
* bcd_in1=00011000 bcd_in2=00100010 cout=0 sum=01000000
* bcd_in1=00011000 bcd_in2=00100011 cout=0 sum=01000001
* bcd_in1=00011000 bcd_in2=00100100 cout=0 sum=01000010
* bcd_in1=00011000 bcd_in2=00100101 cout=0 sum=01000011
* bcd_in1=00011000 bcd_in2=00100110 cout=0 sum=01000100
* bcd_in1=00011000 bcd_in2=00100111 cout=0 sum=01000101
* bcd_in1=00011000 bcd_in2=00101000 cout=0 sum=01000110
* bcd_in1=00011000 bcd_in2=00101001 cout=0 sum=01000111
* bcd_in1=00011000 bcd_in2=00110000 cout=0 sum=01001000
* bcd_in1=00011000 bcd_in2=00110001 cout=0 sum=01001001
* bcd_in1=00011000 bcd_in2=00110010 cout=0 sum=01010000
* bcd_in1=00011000 bcd_in2=00110011 cout=0 sum=01010001
* bcd_in1=00011000 bcd_in2=00110100 cout=0 sum=01010010
* bcd_in1=00011000 bcd_in2=00110101 cout=0 sum=01010011
* bcd_in1=00011000 bcd_in2=00110110 cout=0 sum=01010100
* bcd_in1=00011000 bcd_in2=00110111 cout=0 sum=01010101
* bcd_in1=00011000 bcd_in2=00111000 cout=0 sum=01010110
* bcd_in1=00011000 bcd_in2=00111001 cout=0 sum=01010111
* bcd_in1=00011000 bcd_in2=01000000 cout=0 sum=01011000
* bcd_in1=00011000 bcd_in2=01000001 cout=0 sum=01011001
* bcd_in1=00011000 bcd_in2=01000010 cout=0 sum=01100000
* bcd_in1=00011000 bcd_in2=01000011 cout=0 sum=01100001
* bcd_in1=00011000 bcd_in2=01000100 cout=0 sum=01100010
* bcd_in1=00011000 bcd_in2=01000101 cout=0 sum=01100011
* bcd_in1=00011000 bcd_in2=01000110 cout=0 sum=01100100
* bcd_in1=00011000 bcd_in2=01000111 cout=0 sum=01100101
* bcd_in1=00011000 bcd_in2=01001000 cout=0 sum=01100110
* bcd_in1=00011000 bcd_in2=01001001 cout=0 sum=01100111
* bcd_in1=00011000 bcd_in2=01010000 cout=0 sum=01101000
* bcd_in1=00011000 bcd_in2=01010001 cout=0 sum=01101001
* bcd_in1=00011000 bcd_in2=01010010 cout=0 sum=01110000
* bcd_in1=00011000 bcd_in2=01010011 cout=0 sum=01110001
* bcd_in1=00011000 bcd_in2=01010100 cout=0 sum=01110010
* bcd_in1=00011000 bcd_in2=01010101 cout=0 sum=01110011
* bcd_in1=00011000 bcd_in2=01010110 cout=0 sum=01110100
* bcd_in1=00011000 bcd_in2=01010111 cout=0 sum=01110101
* bcd_in1=00011000 bcd_in2=01011000 cout=0 sum=01110110
* bcd_in1=00011000 bcd_in2=01011001 cout=0 sum=01110111
* bcd_in1=00011000 bcd_in2=01100000 cout=0 sum=01111000
* bcd_in1=00011000 bcd_in2=01100001 cout=0 sum=01111001
* bcd_in1=00011000 bcd_in2=01100010 cout=0 sum=10000000
* bcd_in1=00011000 bcd_in2=01100011 cout=0 sum=10000001
* bcd_in1=00011000 bcd_in2=01100100 cout=0 sum=10000010
* bcd_in1=00011000 bcd_in2=01100101 cout=0 sum=10000011
* bcd_in1=00011000 bcd_in2=01100110 cout=0 sum=10000100
* bcd_in1=00011000 bcd_in2=01100111 cout=0 sum=10000101
* bcd_in1=00011000 bcd_in2=01101000 cout=0 sum=10000110
* bcd_in1=00011000 bcd_in2=01101001 cout=0 sum=10000111
* bcd_in1=00011000 bcd_in2=01110000 cout=0 sum=10001000
* bcd_in1=00011000 bcd_in2=01110001 cout=0 sum=10001001
* bcd_in1=00011000 bcd_in2=01110010 cout=0 sum=10010000
* bcd_in1=00011000 bcd_in2=01110011 cout=0 sum=10010001
* bcd_in1=00011000 bcd_in2=01110100 cout=0 sum=10010010
* bcd_in1=00011000 bcd_in2=01110101 cout=0 sum=10010011
* bcd_in1=00011000 bcd_in2=01110110 cout=0 sum=10010100
* bcd_in1=00011000 bcd_in2=01110111 cout=0 sum=10010101
* bcd_in1=00011000 bcd_in2=01111000 cout=0 sum=10010110
* bcd_in1=00011000 bcd_in2=01111001 cout=0 sum=10010111
* bcd_in1=00011000 bcd_in2=10000000 cout=0 sum=10011000
* bcd_in1=00011000 bcd_in2=10000001 cout=0 sum=10011001
* bcd_in1=00011000 bcd_in2=10000010 cout=1 sum=00000000
* bcd_in1=00011000 bcd_in2=10000011 cout=1 sum=00000001
* bcd_in1=00011000 bcd_in2=10000100 cout=1 sum=00000010
* bcd_in1=00011000 bcd_in2=10000101 cout=1 sum=00000011
* bcd_in1=00011000 bcd_in2=10000110 cout=1 sum=00000100
* bcd_in1=00011000 bcd_in2=10000111 cout=1 sum=00000101
* bcd_in1=00011000 bcd_in2=10001000 cout=1 sum=00000110
* bcd_in1=00011000 bcd_in2=10001001 cout=1 sum=00000111
* bcd_in1=00011000 bcd_in2=10010000 cout=1 sum=00001000
* bcd_in1=00011000 bcd_in2=10010001 cout=1 sum=00001001
* bcd_in1=00011000 bcd_in2=10010010 cout=1 sum=00010000
* bcd_in1=00011000 bcd_in2=10010011 cout=1 sum=00010001
* bcd_in1=00011000 bcd_in2=10010100 cout=1 sum=00010010
* bcd_in1=00011000 bcd_in2=10010101 cout=1 sum=00010011
* bcd_in1=00011000 bcd_in2=10010110 cout=1 sum=00010100
* bcd_in1=00011000 bcd_in2=10010111 cout=1 sum=00010101
* bcd_in1=00011000 bcd_in2=10011000 cout=1 sum=00010110
* bcd_in1=00011000 bcd_in2=10011001 cout=1 sum=00010111
* bcd_in1=00011001 bcd_in2=00000000 cout=0 sum=00011001
* bcd_in1=00011001 bcd_in2=00000001 cout=0 sum=00100000
* bcd_in1=00011001 bcd_in2=00000010 cout=0 sum=00100001
* bcd_in1=00011001 bcd_in2=00000011 cout=0 sum=00100010
* bcd_in1=00011001 bcd_in2=00000100 cout=0 sum=00100011
* bcd_in1=00011001 bcd_in2=00000101 cout=0 sum=00100100
* bcd_in1=00011001 bcd_in2=00000110 cout=0 sum=00100101
* bcd_in1=00011001 bcd_in2=00000111 cout=0 sum=00100110
* bcd_in1=00011001 bcd_in2=00001000 cout=0 sum=00100111
* bcd_in1=00011001 bcd_in2=00001001 cout=0 sum=00101000
* bcd_in1=00011001 bcd_in2=00010000 cout=0 sum=00101001
* bcd_in1=00011001 bcd_in2=00010001 cout=0 sum=00110000
* bcd_in1=00011001 bcd_in2=00010010 cout=0 sum=00110001
* bcd_in1=00011001 bcd_in2=00010011 cout=0 sum=00110010
* bcd_in1=00011001 bcd_in2=00010100 cout=0 sum=00110011
* bcd_in1=00011001 bcd_in2=00010101 cout=0 sum=00110100
* bcd_in1=00011001 bcd_in2=00010110 cout=0 sum=00110101
* bcd_in1=00011001 bcd_in2=00010111 cout=0 sum=00110110
* bcd_in1=00011001 bcd_in2=00011000 cout=0 sum=00110111
* bcd_in1=00011001 bcd_in2=00011001 cout=0 sum=00111000
* bcd_in1=00011001 bcd_in2=00100000 cout=0 sum=00111001
* bcd_in1=00011001 bcd_in2=00100001 cout=0 sum=01000000
* bcd_in1=00011001 bcd_in2=00100010 cout=0 sum=01000001
* bcd_in1=00011001 bcd_in2=00100011 cout=0 sum=01000010
* bcd_in1=00011001 bcd_in2=00100100 cout=0 sum=01000011
* bcd_in1=00011001 bcd_in2=00100101 cout=0 sum=01000100
* bcd_in1=00011001 bcd_in2=00100110 cout=0 sum=01000101
* bcd_in1=00011001 bcd_in2=00100111 cout=0 sum=01000110
* bcd_in1=00011001 bcd_in2=00101000 cout=0 sum=01000111
* bcd_in1=00011001 bcd_in2=00101001 cout=0 sum=01001000
* bcd_in1=00011001 bcd_in2=00110000 cout=0 sum=01001001
* bcd_in1=00011001 bcd_in2=00110001 cout=0 sum=01010000
* bcd_in1=00011001 bcd_in2=00110010 cout=0 sum=01010001
* bcd_in1=00011001 bcd_in2=00110011 cout=0 sum=01010010
* bcd_in1=00011001 bcd_in2=00110100 cout=0 sum=01010011
* bcd_in1=00011001 bcd_in2=00110101 cout=0 sum=01010100
* bcd_in1=00011001 bcd_in2=00110110 cout=0 sum=01010101
* bcd_in1=00011001 bcd_in2=00110111 cout=0 sum=01010110
* bcd_in1=00011001 bcd_in2=00111000 cout=0 sum=01010111
* bcd_in1=00011001 bcd_in2=00111001 cout=0 sum=01011000
* bcd_in1=00011001 bcd_in2=01000000 cout=0 sum=01011001
* bcd_in1=00011001 bcd_in2=01000001 cout=0 sum=01100000
* bcd_in1=00011001 bcd_in2=01000010 cout=0 sum=01100001
* bcd_in1=00011001 bcd_in2=01000011 cout=0 sum=01100010
* bcd_in1=00011001 bcd_in2=01000100 cout=0 sum=01100011
* bcd_in1=00011001 bcd_in2=01000101 cout=0 sum=01100100
* bcd_in1=00011001 bcd_in2=01000110 cout=0 sum=01100101
* bcd_in1=00011001 bcd_in2=01000111 cout=0 sum=01100110
* bcd_in1=00011001 bcd_in2=01001000 cout=0 sum=01100111
* bcd_in1=00011001 bcd_in2=01001001 cout=0 sum=01101000
* bcd_in1=00011001 bcd_in2=01010000 cout=0 sum=01101001
* bcd_in1=00011001 bcd_in2=01010001 cout=0 sum=01110000
* bcd_in1=00011001 bcd_in2=01010010 cout=0 sum=01110001
* bcd_in1=00011001 bcd_in2=01010011 cout=0 sum=01110010
* bcd_in1=00011001 bcd_in2=01010100 cout=0 sum=01110011
* bcd_in1=00011001 bcd_in2=01010101 cout=0 sum=01110100
* bcd_in1=00011001 bcd_in2=01010110 cout=0 sum=01110101
* bcd_in1=00011001 bcd_in2=01010111 cout=0 sum=01110110
* bcd_in1=00011001 bcd_in2=01011000 cout=0 sum=01110111
* bcd_in1=00011001 bcd_in2=01011001 cout=0 sum=01111000
* bcd_in1=00011001 bcd_in2=01100000 cout=0 sum=01111001
* bcd_in1=00011001 bcd_in2=01100001 cout=0 sum=10000000
* bcd_in1=00011001 bcd_in2=01100010 cout=0 sum=10000001
* bcd_in1=00011001 bcd_in2=01100011 cout=0 sum=10000010
* bcd_in1=00011001 bcd_in2=01100100 cout=0 sum=10000011
* bcd_in1=00011001 bcd_in2=01100101 cout=0 sum=10000100
* bcd_in1=00011001 bcd_in2=01100110 cout=0 sum=10000101
* bcd_in1=00011001 bcd_in2=01100111 cout=0 sum=10000110
* bcd_in1=00011001 bcd_in2=01101000 cout=0 sum=10000111
* bcd_in1=00011001 bcd_in2=01101001 cout=0 sum=10001000
* bcd_in1=00011001 bcd_in2=01110000 cout=0 sum=10001001
* bcd_in1=00011001 bcd_in2=01110001 cout=0 sum=10010000
* bcd_in1=00011001 bcd_in2=01110010 cout=0 sum=10010001
* bcd_in1=00011001 bcd_in2=01110011 cout=0 sum=10010010
* bcd_in1=00011001 bcd_in2=01110100 cout=0 sum=10010011
* bcd_in1=00011001 bcd_in2=01110101 cout=0 sum=10010100
* bcd_in1=00011001 bcd_in2=01110110 cout=0 sum=10010101
* bcd_in1=00011001 bcd_in2=01110111 cout=0 sum=10010110
* bcd_in1=00011001 bcd_in2=01111000 cout=0 sum=10010111
* bcd_in1=00011001 bcd_in2=01111001 cout=0 sum=10011000
* bcd_in1=00011001 bcd_in2=10000000 cout=0 sum=10011001
* bcd_in1=00011001 bcd_in2=10000001 cout=1 sum=00000000
* bcd_in1=00011001 bcd_in2=10000010 cout=1 sum=00000001
* bcd_in1=00011001 bcd_in2=10000011 cout=1 sum=00000010
* bcd_in1=00011001 bcd_in2=10000100 cout=1 sum=00000011
* bcd_in1=00011001 bcd_in2=10000101 cout=1 sum=00000100
* bcd_in1=00011001 bcd_in2=10000110 cout=1 sum=00000101
* bcd_in1=00011001 bcd_in2=10000111 cout=1 sum=00000110
* bcd_in1=00011001 bcd_in2=10001000 cout=1 sum=00000111
* bcd_in1=00011001 bcd_in2=10001001 cout=1 sum=00001000
* bcd_in1=00011001 bcd_in2=10010000 cout=1 sum=00001001
* bcd_in1=00011001 bcd_in2=10010001 cout=1 sum=00010000
* bcd_in1=00011001 bcd_in2=10010010 cout=1 sum=00010001
* bcd_in1=00011001 bcd_in2=10010011 cout=1 sum=00010010
* bcd_in1=00011001 bcd_in2=10010100 cout=1 sum=00010011
* bcd_in1=00011001 bcd_in2=10010101 cout=1 sum=00010100
* bcd_in1=00011001 bcd_in2=10010110 cout=1 sum=00010101
* bcd_in1=00011001 bcd_in2=10010111 cout=1 sum=00010110
* bcd_in1=00011001 bcd_in2=10011000 cout=1 sum=00010111
* bcd_in1=00011001 bcd_in2=10011001 cout=1 sum=00011000
* bcd_in1=00100000 bcd_in2=00000000 cout=0 sum=00100000
* bcd_in1=00100000 bcd_in2=00000001 cout=0 sum=00100001
* bcd_in1=00100000 bcd_in2=00000010 cout=0 sum=00100010
* bcd_in1=00100000 bcd_in2=00000011 cout=0 sum=00100011
* bcd_in1=00100000 bcd_in2=00000100 cout=0 sum=00100100
* bcd_in1=00100000 bcd_in2=00000101 cout=0 sum=00100101
* bcd_in1=00100000 bcd_in2=00000110 cout=0 sum=00100110
* bcd_in1=00100000 bcd_in2=00000111 cout=0 sum=00100111
* bcd_in1=00100000 bcd_in2=00001000 cout=0 sum=00101000
* bcd_in1=00100000 bcd_in2=00001001 cout=0 sum=00101001
* bcd_in1=00100000 bcd_in2=00010000 cout=0 sum=00110000
* bcd_in1=00100000 bcd_in2=00010001 cout=0 sum=00110001
* bcd_in1=00100000 bcd_in2=00010010 cout=0 sum=00110010
* bcd_in1=00100000 bcd_in2=00010011 cout=0 sum=00110011
* bcd_in1=00100000 bcd_in2=00010100 cout=0 sum=00110100
* bcd_in1=00100000 bcd_in2=00010101 cout=0 sum=00110101
* bcd_in1=00100000 bcd_in2=00010110 cout=0 sum=00110110
* bcd_in1=00100000 bcd_in2=00010111 cout=0 sum=00110111
* bcd_in1=00100000 bcd_in2=00011000 cout=0 sum=00111000
* bcd_in1=00100000 bcd_in2=00011001 cout=0 sum=00111001
* bcd_in1=00100000 bcd_in2=00100000 cout=0 sum=01000000
* bcd_in1=00100000 bcd_in2=00100001 cout=0 sum=01000001
* bcd_in1=00100000 bcd_in2=00100010 cout=0 sum=01000010
* bcd_in1=00100000 bcd_in2=00100011 cout=0 sum=01000011
* bcd_in1=00100000 bcd_in2=00100100 cout=0 sum=01000100
* bcd_in1=00100000 bcd_in2=00100101 cout=0 sum=01000101
* bcd_in1=00100000 bcd_in2=00100110 cout=0 sum=01000110
* bcd_in1=00100000 bcd_in2=00100111 cout=0 sum=01000111
* bcd_in1=00100000 bcd_in2=00101000 cout=0 sum=01001000
* bcd_in1=00100000 bcd_in2=00101001 cout=0 sum=01001001
* bcd_in1=00100000 bcd_in2=00110000 cout=0 sum=01010000
* bcd_in1=00100000 bcd_in2=00110001 cout=0 sum=01010001
* bcd_in1=00100000 bcd_in2=00110010 cout=0 sum=01010010
* bcd_in1=00100000 bcd_in2=00110011 cout=0 sum=01010011
* bcd_in1=00100000 bcd_in2=00110100 cout=0 sum=01010100
* bcd_in1=00100000 bcd_in2=00110101 cout=0 sum=01010101
* bcd_in1=00100000 bcd_in2=00110110 cout=0 sum=01010110
* bcd_in1=00100000 bcd_in2=00110111 cout=0 sum=01010111
* bcd_in1=00100000 bcd_in2=00111000 cout=0 sum=01011000
* bcd_in1=00100000 bcd_in2=00111001 cout=0 sum=01011001
* bcd_in1=00100000 bcd_in2=01000000 cout=0 sum=01100000
* bcd_in1=00100000 bcd_in2=01000001 cout=0 sum=01100001
* bcd_in1=00100000 bcd_in2=01000010 cout=0 sum=01100010
* bcd_in1=00100000 bcd_in2=01000011 cout=0 sum=01100011
* bcd_in1=00100000 bcd_in2=01000100 cout=0 sum=01100100
* bcd_in1=00100000 bcd_in2=01000101 cout=0 sum=01100101
* bcd_in1=00100000 bcd_in2=01000110 cout=0 sum=01100110
* bcd_in1=00100000 bcd_in2=01000111 cout=0 sum=01100111
* bcd_in1=00100000 bcd_in2=01001000 cout=0 sum=01101000
* bcd_in1=00100000 bcd_in2=01001001 cout=0 sum=01101001
* bcd_in1=00100000 bcd_in2=01010000 cout=0 sum=01110000
* bcd_in1=00100000 bcd_in2=01010001 cout=0 sum=01110001
* bcd_in1=00100000 bcd_in2=01010010 cout=0 sum=01110010
* bcd_in1=00100000 bcd_in2=01010011 cout=0 sum=01110011
* bcd_in1=00100000 bcd_in2=01010100 cout=0 sum=01110100
* bcd_in1=00100000 bcd_in2=01010101 cout=0 sum=01110101
* bcd_in1=00100000 bcd_in2=01010110 cout=0 sum=01110110
* bcd_in1=00100000 bcd_in2=01010111 cout=0 sum=01110111
* bcd_in1=00100000 bcd_in2=01011000 cout=0 sum=01111000
* bcd_in1=00100000 bcd_in2=01011001 cout=0 sum=01111001
* bcd_in1=00100000 bcd_in2=01100000 cout=0 sum=10000000
* bcd_in1=00100000 bcd_in2=01100001 cout=0 sum=10000001
* bcd_in1=00100000 bcd_in2=01100010 cout=0 sum=10000010
* bcd_in1=00100000 bcd_in2=01100011 cout=0 sum=10000011
* bcd_in1=00100000 bcd_in2=01100100 cout=0 sum=10000100
* bcd_in1=00100000 bcd_in2=01100101 cout=0 sum=10000101
* bcd_in1=00100000 bcd_in2=01100110 cout=0 sum=10000110
* bcd_in1=00100000 bcd_in2=01100111 cout=0 sum=10000111
* bcd_in1=00100000 bcd_in2=01101000 cout=0 sum=10001000
* bcd_in1=00100000 bcd_in2=01101001 cout=0 sum=10001001
* bcd_in1=00100000 bcd_in2=01110000 cout=0 sum=10010000
* bcd_in1=00100000 bcd_in2=01110001 cout=0 sum=10010001
* bcd_in1=00100000 bcd_in2=01110010 cout=0 sum=10010010
* bcd_in1=00100000 bcd_in2=01110011 cout=0 sum=10010011
* bcd_in1=00100000 bcd_in2=01110100 cout=0 sum=10010100
* bcd_in1=00100000 bcd_in2=01110101 cout=0 sum=10010101
* bcd_in1=00100000 bcd_in2=01110110 cout=0 sum=10010110
* bcd_in1=00100000 bcd_in2=01110111 cout=0 sum=10010111
* bcd_in1=00100000 bcd_in2=01111000 cout=0 sum=10011000
* bcd_in1=00100000 bcd_in2=01111001 cout=0 sum=10011001
* bcd_in1=00100000 bcd_in2=10000000 cout=1 sum=00000000
* bcd_in1=00100000 bcd_in2=10000001 cout=1 sum=00000001
* bcd_in1=00100000 bcd_in2=10000010 cout=1 sum=00000010
* bcd_in1=00100000 bcd_in2=10000011 cout=1 sum=00000011
* bcd_in1=00100000 bcd_in2=10000100 cout=1 sum=00000100
* bcd_in1=00100000 bcd_in2=10000101 cout=1 sum=00000101
* bcd_in1=00100000 bcd_in2=10000110 cout=1 sum=00000110
* bcd_in1=00100000 bcd_in2=10000111 cout=1 sum=00000111
* bcd_in1=00100000 bcd_in2=10001000 cout=1 sum=00001000
* bcd_in1=00100000 bcd_in2=10001001 cout=1 sum=00001001
* bcd_in1=00100000 bcd_in2=10010000 cout=1 sum=00010000
* bcd_in1=00100000 bcd_in2=10010001 cout=1 sum=00010001
* bcd_in1=00100000 bcd_in2=10010010 cout=1 sum=00010010
* bcd_in1=00100000 bcd_in2=10010011 cout=1 sum=00010011
* bcd_in1=00100000 bcd_in2=10010100 cout=1 sum=00010100
* bcd_in1=00100000 bcd_in2=10010101 cout=1 sum=00010101
* bcd_in1=00100000 bcd_in2=10010110 cout=1 sum=00010110
* bcd_in1=00100000 bcd_in2=10010111 cout=1 sum=00010111
* bcd_in1=00100000 bcd_in2=10011000 cout=1 sum=00011000
* bcd_in1=00100000 bcd_in2=10011001 cout=1 sum=00011001
* bcd_in1=00100001 bcd_in2=00000000 cout=0 sum=00100001
* bcd_in1=00100001 bcd_in2=00000001 cout=0 sum=00100010
* bcd_in1=00100001 bcd_in2=00000010 cout=0 sum=00100011
* bcd_in1=00100001 bcd_in2=00000011 cout=0 sum=00100100
* bcd_in1=00100001 bcd_in2=00000100 cout=0 sum=00100101
* bcd_in1=00100001 bcd_in2=00000101 cout=0 sum=00100110
* bcd_in1=00100001 bcd_in2=00000110 cout=0 sum=00100111
* bcd_in1=00100001 bcd_in2=00000111 cout=0 sum=00101000
* bcd_in1=00100001 bcd_in2=00001000 cout=0 sum=00101001
* bcd_in1=00100001 bcd_in2=00001001 cout=0 sum=00110000
* bcd_in1=00100001 bcd_in2=00010000 cout=0 sum=00110001
* bcd_in1=00100001 bcd_in2=00010001 cout=0 sum=00110010
* bcd_in1=00100001 bcd_in2=00010010 cout=0 sum=00110011
* bcd_in1=00100001 bcd_in2=00010011 cout=0 sum=00110100
* bcd_in1=00100001 bcd_in2=00010100 cout=0 sum=00110101
* bcd_in1=00100001 bcd_in2=00010101 cout=0 sum=00110110
* bcd_in1=00100001 bcd_in2=00010110 cout=0 sum=00110111
* bcd_in1=00100001 bcd_in2=00010111 cout=0 sum=00111000
* bcd_in1=00100001 bcd_in2=00011000 cout=0 sum=00111001
* bcd_in1=00100001 bcd_in2=00011001 cout=0 sum=01000000
* bcd_in1=00100001 bcd_in2=00100000 cout=0 sum=01000001
* bcd_in1=00100001 bcd_in2=00100001 cout=0 sum=01000010
* bcd_in1=00100001 bcd_in2=00100010 cout=0 sum=01000011
* bcd_in1=00100001 bcd_in2=00100011 cout=0 sum=01000100
* bcd_in1=00100001 bcd_in2=00100100 cout=0 sum=01000101
* bcd_in1=00100001 bcd_in2=00100101 cout=0 sum=01000110
* bcd_in1=00100001 bcd_in2=00100110 cout=0 sum=01000111
* bcd_in1=00100001 bcd_in2=00100111 cout=0 sum=01001000
* bcd_in1=00100001 bcd_in2=00101000 cout=0 sum=01001001
* bcd_in1=00100001 bcd_in2=00101001 cout=0 sum=01010000
* bcd_in1=00100001 bcd_in2=00110000 cout=0 sum=01010001
* bcd_in1=00100001 bcd_in2=00110001 cout=0 sum=01010010
* bcd_in1=00100001 bcd_in2=00110010 cout=0 sum=01010011
* bcd_in1=00100001 bcd_in2=00110011 cout=0 sum=01010100
* bcd_in1=00100001 bcd_in2=00110100 cout=0 sum=01010101
* bcd_in1=00100001 bcd_in2=00110101 cout=0 sum=01010110
* bcd_in1=00100001 bcd_in2=00110110 cout=0 sum=01010111
* bcd_in1=00100001 bcd_in2=00110111 cout=0 sum=01011000
* bcd_in1=00100001 bcd_in2=00111000 cout=0 sum=01011001
* bcd_in1=00100001 bcd_in2=00111001 cout=0 sum=01100000
* bcd_in1=00100001 bcd_in2=01000000 cout=0 sum=01100001
* bcd_in1=00100001 bcd_in2=01000001 cout=0 sum=01100010
* bcd_in1=00100001 bcd_in2=01000010 cout=0 sum=01100011
* bcd_in1=00100001 bcd_in2=01000011 cout=0 sum=01100100
* bcd_in1=00100001 bcd_in2=01000100 cout=0 sum=01100101
* bcd_in1=00100001 bcd_in2=01000101 cout=0 sum=01100110
* bcd_in1=00100001 bcd_in2=01000110 cout=0 sum=01100111
* bcd_in1=00100001 bcd_in2=01000111 cout=0 sum=01101000
* bcd_in1=00100001 bcd_in2=01001000 cout=0 sum=01101001
* bcd_in1=00100001 bcd_in2=01001001 cout=0 sum=01110000
* bcd_in1=00100001 bcd_in2=01010000 cout=0 sum=01110001
* bcd_in1=00100001 bcd_in2=01010001 cout=0 sum=01110010
* bcd_in1=00100001 bcd_in2=01010010 cout=0 sum=01110011
* bcd_in1=00100001 bcd_in2=01010011 cout=0 sum=01110100
* bcd_in1=00100001 bcd_in2=01010100 cout=0 sum=01110101
* bcd_in1=00100001 bcd_in2=01010101 cout=0 sum=01110110
* bcd_in1=00100001 bcd_in2=01010110 cout=0 sum=01110111
* bcd_in1=00100001 bcd_in2=01010111 cout=0 sum=01111000
* bcd_in1=00100001 bcd_in2=01011000 cout=0 sum=01111001
* bcd_in1=00100001 bcd_in2=01011001 cout=0 sum=10000000
* bcd_in1=00100001 bcd_in2=01100000 cout=0 sum=10000001
* bcd_in1=00100001 bcd_in2=01100001 cout=0 sum=10000010
* bcd_in1=00100001 bcd_in2=01100010 cout=0 sum=10000011
* bcd_in1=00100001 bcd_in2=01100011 cout=0 sum=10000100
* bcd_in1=00100001 bcd_in2=01100100 cout=0 sum=10000101
* bcd_in1=00100001 bcd_in2=01100101 cout=0 sum=10000110
* bcd_in1=00100001 bcd_in2=01100110 cout=0 sum=10000111
* bcd_in1=00100001 bcd_in2=01100111 cout=0 sum=10001000
* bcd_in1=00100001 bcd_in2=01101000 cout=0 sum=10001001
* bcd_in1=00100001 bcd_in2=01101001 cout=0 sum=10010000
* bcd_in1=00100001 bcd_in2=01110000 cout=0 sum=10010001
* bcd_in1=00100001 bcd_in2=01110001 cout=0 sum=10010010
* bcd_in1=00100001 bcd_in2=01110010 cout=0 sum=10010011
* bcd_in1=00100001 bcd_in2=01110011 cout=0 sum=10010100
* bcd_in1=00100001 bcd_in2=01110100 cout=0 sum=10010101
* bcd_in1=00100001 bcd_in2=01110101 cout=0 sum=10010110
* bcd_in1=00100001 bcd_in2=01110110 cout=0 sum=10010111
* bcd_in1=00100001 bcd_in2=01110111 cout=0 sum=10011000
* bcd_in1=00100001 bcd_in2=01111000 cout=0 sum=10011001
* bcd_in1=00100001 bcd_in2=01111001 cout=1 sum=00000000
* bcd_in1=00100001 bcd_in2=10000000 cout=1 sum=00000001
* bcd_in1=00100001 bcd_in2=10000001 cout=1 sum=00000010
* bcd_in1=00100001 bcd_in2=10000010 cout=1 sum=00000011
* bcd_in1=00100001 bcd_in2=10000011 cout=1 sum=00000100
* bcd_in1=00100001 bcd_in2=10000100 cout=1 sum=00000101
* bcd_in1=00100001 bcd_in2=10000101 cout=1 sum=00000110
* bcd_in1=00100001 bcd_in2=10000110 cout=1 sum=00000111
* bcd_in1=00100001 bcd_in2=10000111 cout=1 sum=00001000
* bcd_in1=00100001 bcd_in2=10001000 cout=1 sum=00001001
* bcd_in1=00100001 bcd_in2=10001001 cout=1 sum=00010000
* bcd_in1=00100001 bcd_in2=10010000 cout=1 sum=00010001
* bcd_in1=00100001 bcd_in2=10010001 cout=1 sum=00010010
* bcd_in1=00100001 bcd_in2=10010010 cout=1 sum=00010011
* bcd_in1=00100001 bcd_in2=10010011 cout=1 sum=00010100
* bcd_in1=00100001 bcd_in2=10010100 cout=1 sum=00010101
* bcd_in1=00100001 bcd_in2=10010101 cout=1 sum=00010110
* bcd_in1=00100001 bcd_in2=10010110 cout=1 sum=00010111
* bcd_in1=00100001 bcd_in2=10010111 cout=1 sum=00011000
* bcd_in1=00100001 bcd_in2=10011000 cout=1 sum=00011001
* bcd_in1=00100001 bcd_in2=10011001 cout=1 sum=00100000
* bcd_in1=00100010 bcd_in2=00000000 cout=0 sum=00100010
* bcd_in1=00100010 bcd_in2=00000001 cout=0 sum=00100011
* bcd_in1=00100010 bcd_in2=00000010 cout=0 sum=00100100
* bcd_in1=00100010 bcd_in2=00000011 cout=0 sum=00100101
* bcd_in1=00100010 bcd_in2=00000100 cout=0 sum=00100110
* bcd_in1=00100010 bcd_in2=00000101 cout=0 sum=00100111
* bcd_in1=00100010 bcd_in2=00000110 cout=0 sum=00101000
* bcd_in1=00100010 bcd_in2=00000111 cout=0 sum=00101001
* bcd_in1=00100010 bcd_in2=00001000 cout=0 sum=00110000
* bcd_in1=00100010 bcd_in2=00001001 cout=0 sum=00110001
* bcd_in1=00100010 bcd_in2=00010000 cout=0 sum=00110010
* bcd_in1=00100010 bcd_in2=00010001 cout=0 sum=00110011
* bcd_in1=00100010 bcd_in2=00010010 cout=0 sum=00110100
* bcd_in1=00100010 bcd_in2=00010011 cout=0 sum=00110101
* bcd_in1=00100010 bcd_in2=00010100 cout=0 sum=00110110
* bcd_in1=00100010 bcd_in2=00010101 cout=0 sum=00110111
* bcd_in1=00100010 bcd_in2=00010110 cout=0 sum=00111000
* bcd_in1=00100010 bcd_in2=00010111 cout=0 sum=00111001
* bcd_in1=00100010 bcd_in2=00011000 cout=0 sum=01000000
* bcd_in1=00100010 bcd_in2=00011001 cout=0 sum=01000001
* bcd_in1=00100010 bcd_in2=00100000 cout=0 sum=01000010
* bcd_in1=00100010 bcd_in2=00100001 cout=0 sum=01000011
* bcd_in1=00100010 bcd_in2=00100010 cout=0 sum=01000100
* bcd_in1=00100010 bcd_in2=00100011 cout=0 sum=01000101
* bcd_in1=00100010 bcd_in2=00100100 cout=0 sum=01000110
* bcd_in1=00100010 bcd_in2=00100101 cout=0 sum=01000111
* bcd_in1=00100010 bcd_in2=00100110 cout=0 sum=01001000
* bcd_in1=00100010 bcd_in2=00100111 cout=0 sum=01001001
* bcd_in1=00100010 bcd_in2=00101000 cout=0 sum=01010000
* bcd_in1=00100010 bcd_in2=00101001 cout=0 sum=01010001
* bcd_in1=00100010 bcd_in2=00110000 cout=0 sum=01010010
* bcd_in1=00100010 bcd_in2=00110001 cout=0 sum=01010011
* bcd_in1=00100010 bcd_in2=00110010 cout=0 sum=01010100
* bcd_in1=00100010 bcd_in2=00110011 cout=0 sum=01010101
* bcd_in1=00100010 bcd_in2=00110100 cout=0 sum=01010110
* bcd_in1=00100010 bcd_in2=00110101 cout=0 sum=01010111
* bcd_in1=00100010 bcd_in2=00110110 cout=0 sum=01011000
* bcd_in1=00100010 bcd_in2=00110111 cout=0 sum=01011001
* bcd_in1=00100010 bcd_in2=00111000 cout=0 sum=01100000
* bcd_in1=00100010 bcd_in2=00111001 cout=0 sum=01100001
* bcd_in1=00100010 bcd_in2=01000000 cout=0 sum=01100010
* bcd_in1=00100010 bcd_in2=01000001 cout=0 sum=01100011
* bcd_in1=00100010 bcd_in2=01000010 cout=0 sum=01100100
* bcd_in1=00100010 bcd_in2=01000011 cout=0 sum=01100101
* bcd_in1=00100010 bcd_in2=01000100 cout=0 sum=01100110
* bcd_in1=00100010 bcd_in2=01000101 cout=0 sum=01100111
* bcd_in1=00100010 bcd_in2=01000110 cout=0 sum=01101000
* bcd_in1=00100010 bcd_in2=01000111 cout=0 sum=01101001
* bcd_in1=00100010 bcd_in2=01001000 cout=0 sum=01110000
* bcd_in1=00100010 bcd_in2=01001001 cout=0 sum=01110001
* bcd_in1=00100010 bcd_in2=01010000 cout=0 sum=01110010
* bcd_in1=00100010 bcd_in2=01010001 cout=0 sum=01110011
* bcd_in1=00100010 bcd_in2=01010010 cout=0 sum=01110100
* bcd_in1=00100010 bcd_in2=01010011 cout=0 sum=01110101
* bcd_in1=00100010 bcd_in2=01010100 cout=0 sum=01110110
* bcd_in1=00100010 bcd_in2=01010101 cout=0 sum=01110111
* bcd_in1=00100010 bcd_in2=01010110 cout=0 sum=01111000
* bcd_in1=00100010 bcd_in2=01010111 cout=0 sum=01111001
* bcd_in1=00100010 bcd_in2=01011000 cout=0 sum=10000000
* bcd_in1=00100010 bcd_in2=01011001 cout=0 sum=10000001
* bcd_in1=00100010 bcd_in2=01100000 cout=0 sum=10000010
* bcd_in1=00100010 bcd_in2=01100001 cout=0 sum=10000011
* bcd_in1=00100010 bcd_in2=01100010 cout=0 sum=10000100
* bcd_in1=00100010 bcd_in2=01100011 cout=0 sum=10000101
* bcd_in1=00100010 bcd_in2=01100100 cout=0 sum=10000110
* bcd_in1=00100010 bcd_in2=01100101 cout=0 sum=10000111
* bcd_in1=00100010 bcd_in2=01100110 cout=0 sum=10001000
* bcd_in1=00100010 bcd_in2=01100111 cout=0 sum=10001001
* bcd_in1=00100010 bcd_in2=01101000 cout=0 sum=10010000
* bcd_in1=00100010 bcd_in2=01101001 cout=0 sum=10010001
* bcd_in1=00100010 bcd_in2=01110000 cout=0 sum=10010010
* bcd_in1=00100010 bcd_in2=01110001 cout=0 sum=10010011
* bcd_in1=00100010 bcd_in2=01110010 cout=0 sum=10010100
* bcd_in1=00100010 bcd_in2=01110011 cout=0 sum=10010101
* bcd_in1=00100010 bcd_in2=01110100 cout=0 sum=10010110
* bcd_in1=00100010 bcd_in2=01110101 cout=0 sum=10010111
* bcd_in1=00100010 bcd_in2=01110110 cout=0 sum=10011000
* bcd_in1=00100010 bcd_in2=01110111 cout=0 sum=10011001
* bcd_in1=00100010 bcd_in2=01111000 cout=1 sum=00000000
* bcd_in1=00100010 bcd_in2=01111001 cout=1 sum=00000001
* bcd_in1=00100010 bcd_in2=10000000 cout=1 sum=00000010
* bcd_in1=00100010 bcd_in2=10000001 cout=1 sum=00000011
* bcd_in1=00100010 bcd_in2=10000010 cout=1 sum=00000100
* bcd_in1=00100010 bcd_in2=10000011 cout=1 sum=00000101
* bcd_in1=00100010 bcd_in2=10000100 cout=1 sum=00000110
* bcd_in1=00100010 bcd_in2=10000101 cout=1 sum=00000111
* bcd_in1=00100010 bcd_in2=10000110 cout=1 sum=00001000
* bcd_in1=00100010 bcd_in2=10000111 cout=1 sum=00001001
* bcd_in1=00100010 bcd_in2=10001000 cout=1 sum=00010000
* bcd_in1=00100010 bcd_in2=10001001 cout=1 sum=00010001
* bcd_in1=00100010 bcd_in2=10010000 cout=1 sum=00010010
* bcd_in1=00100010 bcd_in2=10010001 cout=1 sum=00010011
* bcd_in1=00100010 bcd_in2=10010010 cout=1 sum=00010100
* bcd_in1=00100010 bcd_in2=10010011 cout=1 sum=00010101
* bcd_in1=00100010 bcd_in2=10010100 cout=1 sum=00010110
* bcd_in1=00100010 bcd_in2=10010101 cout=1 sum=00010111
* bcd_in1=00100010 bcd_in2=10010110 cout=1 sum=00011000
* bcd_in1=00100010 bcd_in2=10010111 cout=1 sum=00011001
* bcd_in1=00100010 bcd_in2=10011000 cout=1 sum=00100000
* bcd_in1=00100010 bcd_in2=10011001 cout=1 sum=00100001
* bcd_in1=00100011 bcd_in2=00000000 cout=0 sum=00100011
* bcd_in1=00100011 bcd_in2=00000001 cout=0 sum=00100100
* bcd_in1=00100011 bcd_in2=00000010 cout=0 sum=00100101
* bcd_in1=00100011 bcd_in2=00000011 cout=0 sum=00100110
* bcd_in1=00100011 bcd_in2=00000100 cout=0 sum=00100111
* bcd_in1=00100011 bcd_in2=00000101 cout=0 sum=00101000
* bcd_in1=00100011 bcd_in2=00000110 cout=0 sum=00101001
* bcd_in1=00100011 bcd_in2=00000111 cout=0 sum=00110000
* bcd_in1=00100011 bcd_in2=00001000 cout=0 sum=00110001
* bcd_in1=00100011 bcd_in2=00001001 cout=0 sum=00110010
* bcd_in1=00100011 bcd_in2=00010000 cout=0 sum=00110011
* bcd_in1=00100011 bcd_in2=00010001 cout=0 sum=00110100
* bcd_in1=00100011 bcd_in2=00010010 cout=0 sum=00110101
* bcd_in1=00100011 bcd_in2=00010011 cout=0 sum=00110110
* bcd_in1=00100011 bcd_in2=00010100 cout=0 sum=00110111
* bcd_in1=00100011 bcd_in2=00010101 cout=0 sum=00111000
* bcd_in1=00100011 bcd_in2=00010110 cout=0 sum=00111001
* bcd_in1=00100011 bcd_in2=00010111 cout=0 sum=01000000
* bcd_in1=00100011 bcd_in2=00011000 cout=0 sum=01000001
* bcd_in1=00100011 bcd_in2=00011001 cout=0 sum=01000010
* bcd_in1=00100011 bcd_in2=00100000 cout=0 sum=01000011
* bcd_in1=00100011 bcd_in2=00100001 cout=0 sum=01000100
* bcd_in1=00100011 bcd_in2=00100010 cout=0 sum=01000101
* bcd_in1=00100011 bcd_in2=00100011 cout=0 sum=01000110
* bcd_in1=00100011 bcd_in2=00100100 cout=0 sum=01000111
* bcd_in1=00100011 bcd_in2=00100101 cout=0 sum=01001000
* bcd_in1=00100011 bcd_in2=00100110 cout=0 sum=01001001
* bcd_in1=00100011 bcd_in2=00100111 cout=0 sum=01010000
* bcd_in1=00100011 bcd_in2=00101000 cout=0 sum=01010001
* bcd_in1=00100011 bcd_in2=00101001 cout=0 sum=01010010
* bcd_in1=00100011 bcd_in2=00110000 cout=0 sum=01010011
* bcd_in1=00100011 bcd_in2=00110001 cout=0 sum=01010100
* bcd_in1=00100011 bcd_in2=00110010 cout=0 sum=01010101
* bcd_in1=00100011 bcd_in2=00110011 cout=0 sum=01010110
* bcd_in1=00100011 bcd_in2=00110100 cout=0 sum=01010111
* bcd_in1=00100011 bcd_in2=00110101 cout=0 sum=01011000
* bcd_in1=00100011 bcd_in2=00110110 cout=0 sum=01011001
* bcd_in1=00100011 bcd_in2=00110111 cout=0 sum=01100000
* bcd_in1=00100011 bcd_in2=00111000 cout=0 sum=01100001
* bcd_in1=00100011 bcd_in2=00111001 cout=0 sum=01100010
* bcd_in1=00100011 bcd_in2=01000000 cout=0 sum=01100011
* bcd_in1=00100011 bcd_in2=01000001 cout=0 sum=01100100
* bcd_in1=00100011 bcd_in2=01000010 cout=0 sum=01100101
* bcd_in1=00100011 bcd_in2=01000011 cout=0 sum=01100110
* bcd_in1=00100011 bcd_in2=01000100 cout=0 sum=01100111
* bcd_in1=00100011 bcd_in2=01000101 cout=0 sum=01101000
* bcd_in1=00100011 bcd_in2=01000110 cout=0 sum=01101001
* bcd_in1=00100011 bcd_in2=01000111 cout=0 sum=01110000
* bcd_in1=00100011 bcd_in2=01001000 cout=0 sum=01110001
* bcd_in1=00100011 bcd_in2=01001001 cout=0 sum=01110010
* bcd_in1=00100011 bcd_in2=01010000 cout=0 sum=01110011
* bcd_in1=00100011 bcd_in2=01010001 cout=0 sum=01110100
* bcd_in1=00100011 bcd_in2=01010010 cout=0 sum=01110101
* bcd_in1=00100011 bcd_in2=01010011 cout=0 sum=01110110
* bcd_in1=00100011 bcd_in2=01010100 cout=0 sum=01110111
* bcd_in1=00100011 bcd_in2=01010101 cout=0 sum=01111000
* bcd_in1=00100011 bcd_in2=01010110 cout=0 sum=01111001
* bcd_in1=00100011 bcd_in2=01010111 cout=0 sum=10000000
* bcd_in1=00100011 bcd_in2=01011000 cout=0 sum=10000001
* bcd_in1=00100011 bcd_in2=01011001 cout=0 sum=10000010
* bcd_in1=00100011 bcd_in2=01100000 cout=0 sum=10000011
* bcd_in1=00100011 bcd_in2=01100001 cout=0 sum=10000100
* bcd_in1=00100011 bcd_in2=01100010 cout=0 sum=10000101
* bcd_in1=00100011 bcd_in2=01100011 cout=0 sum=10000110
* bcd_in1=00100011 bcd_in2=01100100 cout=0 sum=10000111
* bcd_in1=00100011 bcd_in2=01100101 cout=0 sum=10001000
* bcd_in1=00100011 bcd_in2=01100110 cout=0 sum=10001001
* bcd_in1=00100011 bcd_in2=01100111 cout=0 sum=10010000
* bcd_in1=00100011 bcd_in2=01101000 cout=0 sum=10010001
* bcd_in1=00100011 bcd_in2=01101001 cout=0 sum=10010010
* bcd_in1=00100011 bcd_in2=01110000 cout=0 sum=10010011
* bcd_in1=00100011 bcd_in2=01110001 cout=0 sum=10010100
* bcd_in1=00100011 bcd_in2=01110010 cout=0 sum=10010101
* bcd_in1=00100011 bcd_in2=01110011 cout=0 sum=10010110
* bcd_in1=00100011 bcd_in2=01110100 cout=0 sum=10010111
* bcd_in1=00100011 bcd_in2=01110101 cout=0 sum=10011000
* bcd_in1=00100011 bcd_in2=01110110 cout=0 sum=10011001
* bcd_in1=00100011 bcd_in2=01110111 cout=1 sum=00000000
* bcd_in1=00100011 bcd_in2=01111000 cout=1 sum=00000001
* bcd_in1=00100011 bcd_in2=01111001 cout=1 sum=00000010
* bcd_in1=00100011 bcd_in2=10000000 cout=1 sum=00000011
* bcd_in1=00100011 bcd_in2=10000001 cout=1 sum=00000100
* bcd_in1=00100011 bcd_in2=10000010 cout=1 sum=00000101
* bcd_in1=00100011 bcd_in2=10000011 cout=1 sum=00000110
* bcd_in1=00100011 bcd_in2=10000100 cout=1 sum=00000111
* bcd_in1=00100011 bcd_in2=10000101 cout=1 sum=00001000
* bcd_in1=00100011 bcd_in2=10000110 cout=1 sum=00001001
* bcd_in1=00100011 bcd_in2=10000111 cout=1 sum=00010000
* bcd_in1=00100011 bcd_in2=10001000 cout=1 sum=00010001
* bcd_in1=00100011 bcd_in2=10001001 cout=1 sum=00010010
* bcd_in1=00100011 bcd_in2=10010000 cout=1 sum=00010011
* bcd_in1=00100011 bcd_in2=10010001 cout=1 sum=00010100
* bcd_in1=00100011 bcd_in2=10010010 cout=1 sum=00010101
* bcd_in1=00100011 bcd_in2=10010011 cout=1 sum=00010110
* bcd_in1=00100011 bcd_in2=10010100 cout=1 sum=00010111
* bcd_in1=00100011 bcd_in2=10010101 cout=1 sum=00011000
* bcd_in1=00100011 bcd_in2=10010110 cout=1 sum=00011001
* bcd_in1=00100011 bcd_in2=10010111 cout=1 sum=00100000
* bcd_in1=00100011 bcd_in2=10011000 cout=1 sum=00100001
* bcd_in1=00100011 bcd_in2=10011001 cout=1 sum=00100010
* bcd_in1=00100100 bcd_in2=00000000 cout=0 sum=00100100
* bcd_in1=00100100 bcd_in2=00000001 cout=0 sum=00100101
* bcd_in1=00100100 bcd_in2=00000010 cout=0 sum=00100110
* bcd_in1=00100100 bcd_in2=00000011 cout=0 sum=00100111
* bcd_in1=00100100 bcd_in2=00000100 cout=0 sum=00101000
* bcd_in1=00100100 bcd_in2=00000101 cout=0 sum=00101001
* bcd_in1=00100100 bcd_in2=00000110 cout=0 sum=00110000
* bcd_in1=00100100 bcd_in2=00000111 cout=0 sum=00110001
* bcd_in1=00100100 bcd_in2=00001000 cout=0 sum=00110010
* bcd_in1=00100100 bcd_in2=00001001 cout=0 sum=00110011
* bcd_in1=00100100 bcd_in2=00010000 cout=0 sum=00110100
* bcd_in1=00100100 bcd_in2=00010001 cout=0 sum=00110101
* bcd_in1=00100100 bcd_in2=00010010 cout=0 sum=00110110
* bcd_in1=00100100 bcd_in2=00010011 cout=0 sum=00110111
* bcd_in1=00100100 bcd_in2=00010100 cout=0 sum=00111000
* bcd_in1=00100100 bcd_in2=00010101 cout=0 sum=00111001
* bcd_in1=00100100 bcd_in2=00010110 cout=0 sum=01000000
* bcd_in1=00100100 bcd_in2=00010111 cout=0 sum=01000001
* bcd_in1=00100100 bcd_in2=00011000 cout=0 sum=01000010
* bcd_in1=00100100 bcd_in2=00011001 cout=0 sum=01000011
* bcd_in1=00100100 bcd_in2=00100000 cout=0 sum=01000100
* bcd_in1=00100100 bcd_in2=00100001 cout=0 sum=01000101
* bcd_in1=00100100 bcd_in2=00100010 cout=0 sum=01000110
* bcd_in1=00100100 bcd_in2=00100011 cout=0 sum=01000111
* bcd_in1=00100100 bcd_in2=00100100 cout=0 sum=01001000
* bcd_in1=00100100 bcd_in2=00100101 cout=0 sum=01001001
* bcd_in1=00100100 bcd_in2=00100110 cout=0 sum=01010000
* bcd_in1=00100100 bcd_in2=00100111 cout=0 sum=01010001
* bcd_in1=00100100 bcd_in2=00101000 cout=0 sum=01010010
* bcd_in1=00100100 bcd_in2=00101001 cout=0 sum=01010011
* bcd_in1=00100100 bcd_in2=00110000 cout=0 sum=01010100
* bcd_in1=00100100 bcd_in2=00110001 cout=0 sum=01010101
* bcd_in1=00100100 bcd_in2=00110010 cout=0 sum=01010110
* bcd_in1=00100100 bcd_in2=00110011 cout=0 sum=01010111
* bcd_in1=00100100 bcd_in2=00110100 cout=0 sum=01011000
* bcd_in1=00100100 bcd_in2=00110101 cout=0 sum=01011001
* bcd_in1=00100100 bcd_in2=00110110 cout=0 sum=01100000
* bcd_in1=00100100 bcd_in2=00110111 cout=0 sum=01100001
* bcd_in1=00100100 bcd_in2=00111000 cout=0 sum=01100010
* bcd_in1=00100100 bcd_in2=00111001 cout=0 sum=01100011
* bcd_in1=00100100 bcd_in2=01000000 cout=0 sum=01100100
* bcd_in1=00100100 bcd_in2=01000001 cout=0 sum=01100101
* bcd_in1=00100100 bcd_in2=01000010 cout=0 sum=01100110
* bcd_in1=00100100 bcd_in2=01000011 cout=0 sum=01100111
* bcd_in1=00100100 bcd_in2=01000100 cout=0 sum=01101000
* bcd_in1=00100100 bcd_in2=01000101 cout=0 sum=01101001
* bcd_in1=00100100 bcd_in2=01000110 cout=0 sum=01110000
* bcd_in1=00100100 bcd_in2=01000111 cout=0 sum=01110001
* bcd_in1=00100100 bcd_in2=01001000 cout=0 sum=01110010
* bcd_in1=00100100 bcd_in2=01001001 cout=0 sum=01110011
* bcd_in1=00100100 bcd_in2=01010000 cout=0 sum=01110100
* bcd_in1=00100100 bcd_in2=01010001 cout=0 sum=01110101
* bcd_in1=00100100 bcd_in2=01010010 cout=0 sum=01110110
* bcd_in1=00100100 bcd_in2=01010011 cout=0 sum=01110111
* bcd_in1=00100100 bcd_in2=01010100 cout=0 sum=01111000
* bcd_in1=00100100 bcd_in2=01010101 cout=0 sum=01111001
* bcd_in1=00100100 bcd_in2=01010110 cout=0 sum=10000000
* bcd_in1=00100100 bcd_in2=01010111 cout=0 sum=10000001
* bcd_in1=00100100 bcd_in2=01011000 cout=0 sum=10000010
* bcd_in1=00100100 bcd_in2=01011001 cout=0 sum=10000011
* bcd_in1=00100100 bcd_in2=01100000 cout=0 sum=10000100
* bcd_in1=00100100 bcd_in2=01100001 cout=0 sum=10000101
* bcd_in1=00100100 bcd_in2=01100010 cout=0 sum=10000110
* bcd_in1=00100100 bcd_in2=01100011 cout=0 sum=10000111
* bcd_in1=00100100 bcd_in2=01100100 cout=0 sum=10001000
* bcd_in1=00100100 bcd_in2=01100101 cout=0 sum=10001001
* bcd_in1=00100100 bcd_in2=01100110 cout=0 sum=10010000
* bcd_in1=00100100 bcd_in2=01100111 cout=0 sum=10010001
* bcd_in1=00100100 bcd_in2=01101000 cout=0 sum=10010010
* bcd_in1=00100100 bcd_in2=01101001 cout=0 sum=10010011
* bcd_in1=00100100 bcd_in2=01110000 cout=0 sum=10010100
* bcd_in1=00100100 bcd_in2=01110001 cout=0 sum=10010101
* bcd_in1=00100100 bcd_in2=01110010 cout=0 sum=10010110
* bcd_in1=00100100 bcd_in2=01110011 cout=0 sum=10010111
* bcd_in1=00100100 bcd_in2=01110100 cout=0 sum=10011000
* bcd_in1=00100100 bcd_in2=01110101 cout=0 sum=10011001
* bcd_in1=00100100 bcd_in2=01110110 cout=1 sum=00000000
* bcd_in1=00100100 bcd_in2=01110111 cout=1 sum=00000001
* bcd_in1=00100100 bcd_in2=01111000 cout=1 sum=00000010
* bcd_in1=00100100 bcd_in2=01111001 cout=1 sum=00000011
* bcd_in1=00100100 bcd_in2=10000000 cout=1 sum=00000100
* bcd_in1=00100100 bcd_in2=10000001 cout=1 sum=00000101
* bcd_in1=00100100 bcd_in2=10000010 cout=1 sum=00000110
* bcd_in1=00100100 bcd_in2=10000011 cout=1 sum=00000111
* bcd_in1=00100100 bcd_in2=10000100 cout=1 sum=00001000
* bcd_in1=00100100 bcd_in2=10000101 cout=1 sum=00001001
* bcd_in1=00100100 bcd_in2=10000110 cout=1 sum=00010000
* bcd_in1=00100100 bcd_in2=10000111 cout=1 sum=00010001
* bcd_in1=00100100 bcd_in2=10001000 cout=1 sum=00010010
* bcd_in1=00100100 bcd_in2=10001001 cout=1 sum=00010011
* bcd_in1=00100100 bcd_in2=10010000 cout=1 sum=00010100
* bcd_in1=00100100 bcd_in2=10010001 cout=1 sum=00010101
* bcd_in1=00100100 bcd_in2=10010010 cout=1 sum=00010110
* bcd_in1=00100100 bcd_in2=10010011 cout=1 sum=00010111
* bcd_in1=00100100 bcd_in2=10010100 cout=1 sum=00011000
* bcd_in1=00100100 bcd_in2=10010101 cout=1 sum=00011001
* bcd_in1=00100100 bcd_in2=10010110 cout=1 sum=00100000
* bcd_in1=00100100 bcd_in2=10010111 cout=1 sum=00100001
* bcd_in1=00100100 bcd_in2=10011000 cout=1 sum=00100010
* bcd_in1=00100100 bcd_in2=10011001 cout=1 sum=00100011
* bcd_in1=00100101 bcd_in2=00000000 cout=0 sum=00100101
* bcd_in1=00100101 bcd_in2=00000001 cout=0 sum=00100110
* bcd_in1=00100101 bcd_in2=00000010 cout=0 sum=00100111
* bcd_in1=00100101 bcd_in2=00000011 cout=0 sum=00101000
* bcd_in1=00100101 bcd_in2=00000100 cout=0 sum=00101001
* bcd_in1=00100101 bcd_in2=00000101 cout=0 sum=00110000
* bcd_in1=00100101 bcd_in2=00000110 cout=0 sum=00110001
* bcd_in1=00100101 bcd_in2=00000111 cout=0 sum=00110010
* bcd_in1=00100101 bcd_in2=00001000 cout=0 sum=00110011
* bcd_in1=00100101 bcd_in2=00001001 cout=0 sum=00110100
* bcd_in1=00100101 bcd_in2=00010000 cout=0 sum=00110101
* bcd_in1=00100101 bcd_in2=00010001 cout=0 sum=00110110
* bcd_in1=00100101 bcd_in2=00010010 cout=0 sum=00110111
* bcd_in1=00100101 bcd_in2=00010011 cout=0 sum=00111000
* bcd_in1=00100101 bcd_in2=00010100 cout=0 sum=00111001
* bcd_in1=00100101 bcd_in2=00010101 cout=0 sum=01000000
* bcd_in1=00100101 bcd_in2=00010110 cout=0 sum=01000001
* bcd_in1=00100101 bcd_in2=00010111 cout=0 sum=01000010
* bcd_in1=00100101 bcd_in2=00011000 cout=0 sum=01000011
* bcd_in1=00100101 bcd_in2=00011001 cout=0 sum=01000100
* bcd_in1=00100101 bcd_in2=00100000 cout=0 sum=01000101
* bcd_in1=00100101 bcd_in2=00100001 cout=0 sum=01000110
* bcd_in1=00100101 bcd_in2=00100010 cout=0 sum=01000111
* bcd_in1=00100101 bcd_in2=00100011 cout=0 sum=01001000
* bcd_in1=00100101 bcd_in2=00100100 cout=0 sum=01001001
* bcd_in1=00100101 bcd_in2=00100101 cout=0 sum=01010000
* bcd_in1=00100101 bcd_in2=00100110 cout=0 sum=01010001
* bcd_in1=00100101 bcd_in2=00100111 cout=0 sum=01010010
* bcd_in1=00100101 bcd_in2=00101000 cout=0 sum=01010011
* bcd_in1=00100101 bcd_in2=00101001 cout=0 sum=01010100
* bcd_in1=00100101 bcd_in2=00110000 cout=0 sum=01010101
* bcd_in1=00100101 bcd_in2=00110001 cout=0 sum=01010110
* bcd_in1=00100101 bcd_in2=00110010 cout=0 sum=01010111
* bcd_in1=00100101 bcd_in2=00110011 cout=0 sum=01011000
* bcd_in1=00100101 bcd_in2=00110100 cout=0 sum=01011001
* bcd_in1=00100101 bcd_in2=00110101 cout=0 sum=01100000
* bcd_in1=00100101 bcd_in2=00110110 cout=0 sum=01100001
* bcd_in1=00100101 bcd_in2=00110111 cout=0 sum=01100010
* bcd_in1=00100101 bcd_in2=00111000 cout=0 sum=01100011
* bcd_in1=00100101 bcd_in2=00111001 cout=0 sum=01100100
* bcd_in1=00100101 bcd_in2=01000000 cout=0 sum=01100101
* bcd_in1=00100101 bcd_in2=01000001 cout=0 sum=01100110
* bcd_in1=00100101 bcd_in2=01000010 cout=0 sum=01100111
* bcd_in1=00100101 bcd_in2=01000011 cout=0 sum=01101000
* bcd_in1=00100101 bcd_in2=01000100 cout=0 sum=01101001
* bcd_in1=00100101 bcd_in2=01000101 cout=0 sum=01110000
* bcd_in1=00100101 bcd_in2=01000110 cout=0 sum=01110001
* bcd_in1=00100101 bcd_in2=01000111 cout=0 sum=01110010
* bcd_in1=00100101 bcd_in2=01001000 cout=0 sum=01110011
* bcd_in1=00100101 bcd_in2=01001001 cout=0 sum=01110100
* bcd_in1=00100101 bcd_in2=01010000 cout=0 sum=01110101
* bcd_in1=00100101 bcd_in2=01010001 cout=0 sum=01110110
* bcd_in1=00100101 bcd_in2=01010010 cout=0 sum=01110111
* bcd_in1=00100101 bcd_in2=01010011 cout=0 sum=01111000
* bcd_in1=00100101 bcd_in2=01010100 cout=0 sum=01111001
* bcd_in1=00100101 bcd_in2=01010101 cout=0 sum=10000000
* bcd_in1=00100101 bcd_in2=01010110 cout=0 sum=10000001
* bcd_in1=00100101 bcd_in2=01010111 cout=0 sum=10000010
* bcd_in1=00100101 bcd_in2=01011000 cout=0 sum=10000011
* bcd_in1=00100101 bcd_in2=01011001 cout=0 sum=10000100
* bcd_in1=00100101 bcd_in2=01100000 cout=0 sum=10000101
* bcd_in1=00100101 bcd_in2=01100001 cout=0 sum=10000110
* bcd_in1=00100101 bcd_in2=01100010 cout=0 sum=10000111
* bcd_in1=00100101 bcd_in2=01100011 cout=0 sum=10001000
* bcd_in1=00100101 bcd_in2=01100100 cout=0 sum=10001001
* bcd_in1=00100101 bcd_in2=01100101 cout=0 sum=10010000
* bcd_in1=00100101 bcd_in2=01100110 cout=0 sum=10010001
* bcd_in1=00100101 bcd_in2=01100111 cout=0 sum=10010010
* bcd_in1=00100101 bcd_in2=01101000 cout=0 sum=10010011
* bcd_in1=00100101 bcd_in2=01101001 cout=0 sum=10010100
* bcd_in1=00100101 bcd_in2=01110000 cout=0 sum=10010101
* bcd_in1=00100101 bcd_in2=01110001 cout=0 sum=10010110
* bcd_in1=00100101 bcd_in2=01110010 cout=0 sum=10010111
* bcd_in1=00100101 bcd_in2=01110011 cout=0 sum=10011000
* bcd_in1=00100101 bcd_in2=01110100 cout=0 sum=10011001
* bcd_in1=00100101 bcd_in2=01110101 cout=1 sum=00000000
* bcd_in1=00100101 bcd_in2=01110110 cout=1 sum=00000001
* bcd_in1=00100101 bcd_in2=01110111 cout=1 sum=00000010
* bcd_in1=00100101 bcd_in2=01111000 cout=1 sum=00000011
* bcd_in1=00100101 bcd_in2=01111001 cout=1 sum=00000100
* bcd_in1=00100101 bcd_in2=10000000 cout=1 sum=00000101
* bcd_in1=00100101 bcd_in2=10000001 cout=1 sum=00000110
* bcd_in1=00100101 bcd_in2=10000010 cout=1 sum=00000111
* bcd_in1=00100101 bcd_in2=10000011 cout=1 sum=00001000
* bcd_in1=00100101 bcd_in2=10000100 cout=1 sum=00001001
* bcd_in1=00100101 bcd_in2=10000101 cout=1 sum=00010000
* bcd_in1=00100101 bcd_in2=10000110 cout=1 sum=00010001
* bcd_in1=00100101 bcd_in2=10000111 cout=1 sum=00010010
* bcd_in1=00100101 bcd_in2=10001000 cout=1 sum=00010011
* bcd_in1=00100101 bcd_in2=10001001 cout=1 sum=00010100
* bcd_in1=00100101 bcd_in2=10010000 cout=1 sum=00010101
* bcd_in1=00100101 bcd_in2=10010001 cout=1 sum=00010110
* bcd_in1=00100101 bcd_in2=10010010 cout=1 sum=00010111
* bcd_in1=00100101 bcd_in2=10010011 cout=1 sum=00011000
* bcd_in1=00100101 bcd_in2=10010100 cout=1 sum=00011001
* bcd_in1=00100101 bcd_in2=10010101 cout=1 sum=00100000
* bcd_in1=00100101 bcd_in2=10010110 cout=1 sum=00100001
* bcd_in1=00100101 bcd_in2=10010111 cout=1 sum=00100010
* bcd_in1=00100101 bcd_in2=10011000 cout=1 sum=00100011
* bcd_in1=00100101 bcd_in2=10011001 cout=1 sum=00100100
* bcd_in1=00100110 bcd_in2=00000000 cout=0 sum=00100110
* bcd_in1=00100110 bcd_in2=00000001 cout=0 sum=00100111
* bcd_in1=00100110 bcd_in2=00000010 cout=0 sum=00101000
* bcd_in1=00100110 bcd_in2=00000011 cout=0 sum=00101001
* bcd_in1=00100110 bcd_in2=00000100 cout=0 sum=00110000
* bcd_in1=00100110 bcd_in2=00000101 cout=0 sum=00110001
* bcd_in1=00100110 bcd_in2=00000110 cout=0 sum=00110010
* bcd_in1=00100110 bcd_in2=00000111 cout=0 sum=00110011
* bcd_in1=00100110 bcd_in2=00001000 cout=0 sum=00110100
* bcd_in1=00100110 bcd_in2=00001001 cout=0 sum=00110101
* bcd_in1=00100110 bcd_in2=00010000 cout=0 sum=00110110
* bcd_in1=00100110 bcd_in2=00010001 cout=0 sum=00110111
* bcd_in1=00100110 bcd_in2=00010010 cout=0 sum=00111000
* bcd_in1=00100110 bcd_in2=00010011 cout=0 sum=00111001
* bcd_in1=00100110 bcd_in2=00010100 cout=0 sum=01000000
* bcd_in1=00100110 bcd_in2=00010101 cout=0 sum=01000001
* bcd_in1=00100110 bcd_in2=00010110 cout=0 sum=01000010
* bcd_in1=00100110 bcd_in2=00010111 cout=0 sum=01000011
* bcd_in1=00100110 bcd_in2=00011000 cout=0 sum=01000100
* bcd_in1=00100110 bcd_in2=00011001 cout=0 sum=01000101
* bcd_in1=00100110 bcd_in2=00100000 cout=0 sum=01000110
* bcd_in1=00100110 bcd_in2=00100001 cout=0 sum=01000111
* bcd_in1=00100110 bcd_in2=00100010 cout=0 sum=01001000
* bcd_in1=00100110 bcd_in2=00100011 cout=0 sum=01001001
* bcd_in1=00100110 bcd_in2=00100100 cout=0 sum=01010000
* bcd_in1=00100110 bcd_in2=00100101 cout=0 sum=01010001
* bcd_in1=00100110 bcd_in2=00100110 cout=0 sum=01010010
* bcd_in1=00100110 bcd_in2=00100111 cout=0 sum=01010011
* bcd_in1=00100110 bcd_in2=00101000 cout=0 sum=01010100
* bcd_in1=00100110 bcd_in2=00101001 cout=0 sum=01010101
* bcd_in1=00100110 bcd_in2=00110000 cout=0 sum=01010110
* bcd_in1=00100110 bcd_in2=00110001 cout=0 sum=01010111
* bcd_in1=00100110 bcd_in2=00110010 cout=0 sum=01011000
* bcd_in1=00100110 bcd_in2=00110011 cout=0 sum=01011001
* bcd_in1=00100110 bcd_in2=00110100 cout=0 sum=01100000
* bcd_in1=00100110 bcd_in2=00110101 cout=0 sum=01100001
* bcd_in1=00100110 bcd_in2=00110110 cout=0 sum=01100010
* bcd_in1=00100110 bcd_in2=00110111 cout=0 sum=01100011
* bcd_in1=00100110 bcd_in2=00111000 cout=0 sum=01100100
* bcd_in1=00100110 bcd_in2=00111001 cout=0 sum=01100101
* bcd_in1=00100110 bcd_in2=01000000 cout=0 sum=01100110
* bcd_in1=00100110 bcd_in2=01000001 cout=0 sum=01100111
* bcd_in1=00100110 bcd_in2=01000010 cout=0 sum=01101000
* bcd_in1=00100110 bcd_in2=01000011 cout=0 sum=01101001
* bcd_in1=00100110 bcd_in2=01000100 cout=0 sum=01110000
* bcd_in1=00100110 bcd_in2=01000101 cout=0 sum=01110001
* bcd_in1=00100110 bcd_in2=01000110 cout=0 sum=01110010
* bcd_in1=00100110 bcd_in2=01000111 cout=0 sum=01110011
* bcd_in1=00100110 bcd_in2=01001000 cout=0 sum=01110100
* bcd_in1=00100110 bcd_in2=01001001 cout=0 sum=01110101
* bcd_in1=00100110 bcd_in2=01010000 cout=0 sum=01110110
* bcd_in1=00100110 bcd_in2=01010001 cout=0 sum=01110111
* bcd_in1=00100110 bcd_in2=01010010 cout=0 sum=01111000
* bcd_in1=00100110 bcd_in2=01010011 cout=0 sum=01111001
* bcd_in1=00100110 bcd_in2=01010100 cout=0 sum=10000000
* bcd_in1=00100110 bcd_in2=01010101 cout=0 sum=10000001
* bcd_in1=00100110 bcd_in2=01010110 cout=0 sum=10000010
* bcd_in1=00100110 bcd_in2=01010111 cout=0 sum=10000011
* bcd_in1=00100110 bcd_in2=01011000 cout=0 sum=10000100
* bcd_in1=00100110 bcd_in2=01011001 cout=0 sum=10000101
* bcd_in1=00100110 bcd_in2=01100000 cout=0 sum=10000110
* bcd_in1=00100110 bcd_in2=01100001 cout=0 sum=10000111
* bcd_in1=00100110 bcd_in2=01100010 cout=0 sum=10001000
* bcd_in1=00100110 bcd_in2=01100011 cout=0 sum=10001001
* bcd_in1=00100110 bcd_in2=01100100 cout=0 sum=10010000
* bcd_in1=00100110 bcd_in2=01100101 cout=0 sum=10010001
* bcd_in1=00100110 bcd_in2=01100110 cout=0 sum=10010010
* bcd_in1=00100110 bcd_in2=01100111 cout=0 sum=10010011
* bcd_in1=00100110 bcd_in2=01101000 cout=0 sum=10010100
* bcd_in1=00100110 bcd_in2=01101001 cout=0 sum=10010101
* bcd_in1=00100110 bcd_in2=01110000 cout=0 sum=10010110
* bcd_in1=00100110 bcd_in2=01110001 cout=0 sum=10010111
* bcd_in1=00100110 bcd_in2=01110010 cout=0 sum=10011000
* bcd_in1=00100110 bcd_in2=01110011 cout=0 sum=10011001
* bcd_in1=00100110 bcd_in2=01110100 cout=1 sum=00000000
* bcd_in1=00100110 bcd_in2=01110101 cout=1 sum=00000001
* bcd_in1=00100110 bcd_in2=01110110 cout=1 sum=00000010
* bcd_in1=00100110 bcd_in2=01110111 cout=1 sum=00000011
* bcd_in1=00100110 bcd_in2=01111000 cout=1 sum=00000100
* bcd_in1=00100110 bcd_in2=01111001 cout=1 sum=00000101
* bcd_in1=00100110 bcd_in2=10000000 cout=1 sum=00000110
* bcd_in1=00100110 bcd_in2=10000001 cout=1 sum=00000111
* bcd_in1=00100110 bcd_in2=10000010 cout=1 sum=00001000
* bcd_in1=00100110 bcd_in2=10000011 cout=1 sum=00001001
* bcd_in1=00100110 bcd_in2=10000100 cout=1 sum=00010000
* bcd_in1=00100110 bcd_in2=10000101 cout=1 sum=00010001
* bcd_in1=00100110 bcd_in2=10000110 cout=1 sum=00010010
* bcd_in1=00100110 bcd_in2=10000111 cout=1 sum=00010011
* bcd_in1=00100110 bcd_in2=10001000 cout=1 sum=00010100
* bcd_in1=00100110 bcd_in2=10001001 cout=1 sum=00010101
* bcd_in1=00100110 bcd_in2=10010000 cout=1 sum=00010110
* bcd_in1=00100110 bcd_in2=10010001 cout=1 sum=00010111
* bcd_in1=00100110 bcd_in2=10010010 cout=1 sum=00011000
* bcd_in1=00100110 bcd_in2=10010011 cout=1 sum=00011001
* bcd_in1=00100110 bcd_in2=10010100 cout=1 sum=00100000
* bcd_in1=00100110 bcd_in2=10010101 cout=1 sum=00100001
* bcd_in1=00100110 bcd_in2=10010110 cout=1 sum=00100010
* bcd_in1=00100110 bcd_in2=10010111 cout=1 sum=00100011
* bcd_in1=00100110 bcd_in2=10011000 cout=1 sum=00100100
* bcd_in1=00100110 bcd_in2=10011001 cout=1 sum=00100101
* bcd_in1=00100111 bcd_in2=00000000 cout=0 sum=00100111
* bcd_in1=00100111 bcd_in2=00000001 cout=0 sum=00101000
* bcd_in1=00100111 bcd_in2=00000010 cout=0 sum=00101001
* bcd_in1=00100111 bcd_in2=00000011 cout=0 sum=00110000
* bcd_in1=00100111 bcd_in2=00000100 cout=0 sum=00110001
* bcd_in1=00100111 bcd_in2=00000101 cout=0 sum=00110010
* bcd_in1=00100111 bcd_in2=00000110 cout=0 sum=00110011
* bcd_in1=00100111 bcd_in2=00000111 cout=0 sum=00110100
* bcd_in1=00100111 bcd_in2=00001000 cout=0 sum=00110101
* bcd_in1=00100111 bcd_in2=00001001 cout=0 sum=00110110
* bcd_in1=00100111 bcd_in2=00010000 cout=0 sum=00110111
* bcd_in1=00100111 bcd_in2=00010001 cout=0 sum=00111000
* bcd_in1=00100111 bcd_in2=00010010 cout=0 sum=00111001
* bcd_in1=00100111 bcd_in2=00010011 cout=0 sum=01000000
* bcd_in1=00100111 bcd_in2=00010100 cout=0 sum=01000001
* bcd_in1=00100111 bcd_in2=00010101 cout=0 sum=01000010
* bcd_in1=00100111 bcd_in2=00010110 cout=0 sum=01000011
* bcd_in1=00100111 bcd_in2=00010111 cout=0 sum=01000100
* bcd_in1=00100111 bcd_in2=00011000 cout=0 sum=01000101
* bcd_in1=00100111 bcd_in2=00011001 cout=0 sum=01000110
* bcd_in1=00100111 bcd_in2=00100000 cout=0 sum=01000111
* bcd_in1=00100111 bcd_in2=00100001 cout=0 sum=01001000
* bcd_in1=00100111 bcd_in2=00100010 cout=0 sum=01001001
* bcd_in1=00100111 bcd_in2=00100011 cout=0 sum=01010000
* bcd_in1=00100111 bcd_in2=00100100 cout=0 sum=01010001
* bcd_in1=00100111 bcd_in2=00100101 cout=0 sum=01010010
* bcd_in1=00100111 bcd_in2=00100110 cout=0 sum=01010011
* bcd_in1=00100111 bcd_in2=00100111 cout=0 sum=01010100
* bcd_in1=00100111 bcd_in2=00101000 cout=0 sum=01010101
* bcd_in1=00100111 bcd_in2=00101001 cout=0 sum=01010110
* bcd_in1=00100111 bcd_in2=00110000 cout=0 sum=01010111
* bcd_in1=00100111 bcd_in2=00110001 cout=0 sum=01011000
* bcd_in1=00100111 bcd_in2=00110010 cout=0 sum=01011001
* bcd_in1=00100111 bcd_in2=00110011 cout=0 sum=01100000
* bcd_in1=00100111 bcd_in2=00110100 cout=0 sum=01100001
* bcd_in1=00100111 bcd_in2=00110101 cout=0 sum=01100010
* bcd_in1=00100111 bcd_in2=00110110 cout=0 sum=01100011
* bcd_in1=00100111 bcd_in2=00110111 cout=0 sum=01100100
* bcd_in1=00100111 bcd_in2=00111000 cout=0 sum=01100101
* bcd_in1=00100111 bcd_in2=00111001 cout=0 sum=01100110
* bcd_in1=00100111 bcd_in2=01000000 cout=0 sum=01100111
* bcd_in1=00100111 bcd_in2=01000001 cout=0 sum=01101000
* bcd_in1=00100111 bcd_in2=01000010 cout=0 sum=01101001
* bcd_in1=00100111 bcd_in2=01000011 cout=0 sum=01110000
* bcd_in1=00100111 bcd_in2=01000100 cout=0 sum=01110001
* bcd_in1=00100111 bcd_in2=01000101 cout=0 sum=01110010
* bcd_in1=00100111 bcd_in2=01000110 cout=0 sum=01110011
* bcd_in1=00100111 bcd_in2=01000111 cout=0 sum=01110100
* bcd_in1=00100111 bcd_in2=01001000 cout=0 sum=01110101
* bcd_in1=00100111 bcd_in2=01001001 cout=0 sum=01110110
* bcd_in1=00100111 bcd_in2=01010000 cout=0 sum=01110111
* bcd_in1=00100111 bcd_in2=01010001 cout=0 sum=01111000
* bcd_in1=00100111 bcd_in2=01010010 cout=0 sum=01111001
* bcd_in1=00100111 bcd_in2=01010011 cout=0 sum=10000000
* bcd_in1=00100111 bcd_in2=01010100 cout=0 sum=10000001
* bcd_in1=00100111 bcd_in2=01010101 cout=0 sum=10000010
* bcd_in1=00100111 bcd_in2=01010110 cout=0 sum=10000011
* bcd_in1=00100111 bcd_in2=01010111 cout=0 sum=10000100
* bcd_in1=00100111 bcd_in2=01011000 cout=0 sum=10000101
* bcd_in1=00100111 bcd_in2=01011001 cout=0 sum=10000110
* bcd_in1=00100111 bcd_in2=01100000 cout=0 sum=10000111
* bcd_in1=00100111 bcd_in2=01100001 cout=0 sum=10001000
* bcd_in1=00100111 bcd_in2=01100010 cout=0 sum=10001001
* bcd_in1=00100111 bcd_in2=01100011 cout=0 sum=10010000
* bcd_in1=00100111 bcd_in2=01100100 cout=0 sum=10010001
* bcd_in1=00100111 bcd_in2=01100101 cout=0 sum=10010010
* bcd_in1=00100111 bcd_in2=01100110 cout=0 sum=10010011
* bcd_in1=00100111 bcd_in2=01100111 cout=0 sum=10010100
* bcd_in1=00100111 bcd_in2=01101000 cout=0 sum=10010101
* bcd_in1=00100111 bcd_in2=01101001 cout=0 sum=10010110
* bcd_in1=00100111 bcd_in2=01110000 cout=0 sum=10010111
* bcd_in1=00100111 bcd_in2=01110001 cout=0 sum=10011000
* bcd_in1=00100111 bcd_in2=01110010 cout=0 sum=10011001
* bcd_in1=00100111 bcd_in2=01110011 cout=1 sum=00000000
* bcd_in1=00100111 bcd_in2=01110100 cout=1 sum=00000001
* bcd_in1=00100111 bcd_in2=01110101 cout=1 sum=00000010
* bcd_in1=00100111 bcd_in2=01110110 cout=1 sum=00000011
* bcd_in1=00100111 bcd_in2=01110111 cout=1 sum=00000100
* bcd_in1=00100111 bcd_in2=01111000 cout=1 sum=00000101
* bcd_in1=00100111 bcd_in2=01111001 cout=1 sum=00000110
* bcd_in1=00100111 bcd_in2=10000000 cout=1 sum=00000111
* bcd_in1=00100111 bcd_in2=10000001 cout=1 sum=00001000
* bcd_in1=00100111 bcd_in2=10000010 cout=1 sum=00001001
* bcd_in1=00100111 bcd_in2=10000011 cout=1 sum=00010000
* bcd_in1=00100111 bcd_in2=10000100 cout=1 sum=00010001
* bcd_in1=00100111 bcd_in2=10000101 cout=1 sum=00010010
* bcd_in1=00100111 bcd_in2=10000110 cout=1 sum=00010011
* bcd_in1=00100111 bcd_in2=10000111 cout=1 sum=00010100
* bcd_in1=00100111 bcd_in2=10001000 cout=1 sum=00010101
* bcd_in1=00100111 bcd_in2=10001001 cout=1 sum=00010110
* bcd_in1=00100111 bcd_in2=10010000 cout=1 sum=00010111
* bcd_in1=00100111 bcd_in2=10010001 cout=1 sum=00011000
* bcd_in1=00100111 bcd_in2=10010010 cout=1 sum=00011001
* bcd_in1=00100111 bcd_in2=10010011 cout=1 sum=00100000
* bcd_in1=00100111 bcd_in2=10010100 cout=1 sum=00100001
* bcd_in1=00100111 bcd_in2=10010101 cout=1 sum=00100010
* bcd_in1=00100111 bcd_in2=10010110 cout=1 sum=00100011
* bcd_in1=00100111 bcd_in2=10010111 cout=1 sum=00100100
* bcd_in1=00100111 bcd_in2=10011000 cout=1 sum=00100101
* bcd_in1=00100111 bcd_in2=10011001 cout=1 sum=00100110
* bcd_in1=00101000 bcd_in2=00000000 cout=0 sum=00101000
* bcd_in1=00101000 bcd_in2=00000001 cout=0 sum=00101001
* bcd_in1=00101000 bcd_in2=00000010 cout=0 sum=00110000
* bcd_in1=00101000 bcd_in2=00000011 cout=0 sum=00110001
* bcd_in1=00101000 bcd_in2=00000100 cout=0 sum=00110010
* bcd_in1=00101000 bcd_in2=00000101 cout=0 sum=00110011
* bcd_in1=00101000 bcd_in2=00000110 cout=0 sum=00110100
* bcd_in1=00101000 bcd_in2=00000111 cout=0 sum=00110101
* bcd_in1=00101000 bcd_in2=00001000 cout=0 sum=00110110
* bcd_in1=00101000 bcd_in2=00001001 cout=0 sum=00110111
* bcd_in1=00101000 bcd_in2=00010000 cout=0 sum=00111000
* bcd_in1=00101000 bcd_in2=00010001 cout=0 sum=00111001
* bcd_in1=00101000 bcd_in2=00010010 cout=0 sum=01000000
* bcd_in1=00101000 bcd_in2=00010011 cout=0 sum=01000001
* bcd_in1=00101000 bcd_in2=00010100 cout=0 sum=01000010
* bcd_in1=00101000 bcd_in2=00010101 cout=0 sum=01000011
* bcd_in1=00101000 bcd_in2=00010110 cout=0 sum=01000100
* bcd_in1=00101000 bcd_in2=00010111 cout=0 sum=01000101
* bcd_in1=00101000 bcd_in2=00011000 cout=0 sum=01000110
* bcd_in1=00101000 bcd_in2=00011001 cout=0 sum=01000111
* bcd_in1=00101000 bcd_in2=00100000 cout=0 sum=01001000
* bcd_in1=00101000 bcd_in2=00100001 cout=0 sum=01001001
* bcd_in1=00101000 bcd_in2=00100010 cout=0 sum=01010000
* bcd_in1=00101000 bcd_in2=00100011 cout=0 sum=01010001
* bcd_in1=00101000 bcd_in2=00100100 cout=0 sum=01010010
* bcd_in1=00101000 bcd_in2=00100101 cout=0 sum=01010011
* bcd_in1=00101000 bcd_in2=00100110 cout=0 sum=01010100
* bcd_in1=00101000 bcd_in2=00100111 cout=0 sum=01010101
* bcd_in1=00101000 bcd_in2=00101000 cout=0 sum=01010110
* bcd_in1=00101000 bcd_in2=00101001 cout=0 sum=01010111
* bcd_in1=00101000 bcd_in2=00110000 cout=0 sum=01011000
* bcd_in1=00101000 bcd_in2=00110001 cout=0 sum=01011001
* bcd_in1=00101000 bcd_in2=00110010 cout=0 sum=01100000
* bcd_in1=00101000 bcd_in2=00110011 cout=0 sum=01100001
* bcd_in1=00101000 bcd_in2=00110100 cout=0 sum=01100010
* bcd_in1=00101000 bcd_in2=00110101 cout=0 sum=01100011
* bcd_in1=00101000 bcd_in2=00110110 cout=0 sum=01100100
* bcd_in1=00101000 bcd_in2=00110111 cout=0 sum=01100101
* bcd_in1=00101000 bcd_in2=00111000 cout=0 sum=01100110
* bcd_in1=00101000 bcd_in2=00111001 cout=0 sum=01100111
* bcd_in1=00101000 bcd_in2=01000000 cout=0 sum=01101000
* bcd_in1=00101000 bcd_in2=01000001 cout=0 sum=01101001
* bcd_in1=00101000 bcd_in2=01000010 cout=0 sum=01110000
* bcd_in1=00101000 bcd_in2=01000011 cout=0 sum=01110001
* bcd_in1=00101000 bcd_in2=01000100 cout=0 sum=01110010
* bcd_in1=00101000 bcd_in2=01000101 cout=0 sum=01110011
* bcd_in1=00101000 bcd_in2=01000110 cout=0 sum=01110100
* bcd_in1=00101000 bcd_in2=01000111 cout=0 sum=01110101
* bcd_in1=00101000 bcd_in2=01001000 cout=0 sum=01110110
* bcd_in1=00101000 bcd_in2=01001001 cout=0 sum=01110111
* bcd_in1=00101000 bcd_in2=01010000 cout=0 sum=01111000
* bcd_in1=00101000 bcd_in2=01010001 cout=0 sum=01111001
* bcd_in1=00101000 bcd_in2=01010010 cout=0 sum=10000000
* bcd_in1=00101000 bcd_in2=01010011 cout=0 sum=10000001
* bcd_in1=00101000 bcd_in2=01010100 cout=0 sum=10000010
* bcd_in1=00101000 bcd_in2=01010101 cout=0 sum=10000011
* bcd_in1=00101000 bcd_in2=01010110 cout=0 sum=10000100
* bcd_in1=00101000 bcd_in2=01010111 cout=0 sum=10000101
* bcd_in1=00101000 bcd_in2=01011000 cout=0 sum=10000110
* bcd_in1=00101000 bcd_in2=01011001 cout=0 sum=10000111
* bcd_in1=00101000 bcd_in2=01100000 cout=0 sum=10001000
* bcd_in1=00101000 bcd_in2=01100001 cout=0 sum=10001001
* bcd_in1=00101000 bcd_in2=01100010 cout=0 sum=10010000
* bcd_in1=00101000 bcd_in2=01100011 cout=0 sum=10010001
* bcd_in1=00101000 bcd_in2=01100100 cout=0 sum=10010010
* bcd_in1=00101000 bcd_in2=01100101 cout=0 sum=10010011
* bcd_in1=00101000 bcd_in2=01100110 cout=0 sum=10010100
* bcd_in1=00101000 bcd_in2=01100111 cout=0 sum=10010101
* bcd_in1=00101000 bcd_in2=01101000 cout=0 sum=10010110
* bcd_in1=00101000 bcd_in2=01101001 cout=0 sum=10010111
* bcd_in1=00101000 bcd_in2=01110000 cout=0 sum=10011000
* bcd_in1=00101000 bcd_in2=01110001 cout=0 sum=10011001
* bcd_in1=00101000 bcd_in2=01110010 cout=1 sum=00000000
* bcd_in1=00101000 bcd_in2=01110011 cout=1 sum=00000001
* bcd_in1=00101000 bcd_in2=01110100 cout=1 sum=00000010
* bcd_in1=00101000 bcd_in2=01110101 cout=1 sum=00000011
* bcd_in1=00101000 bcd_in2=01110110 cout=1 sum=00000100
* bcd_in1=00101000 bcd_in2=01110111 cout=1 sum=00000101
* bcd_in1=00101000 bcd_in2=01111000 cout=1 sum=00000110
* bcd_in1=00101000 bcd_in2=01111001 cout=1 sum=00000111
* bcd_in1=00101000 bcd_in2=10000000 cout=1 sum=00001000
* bcd_in1=00101000 bcd_in2=10000001 cout=1 sum=00001001
* bcd_in1=00101000 bcd_in2=10000010 cout=1 sum=00010000
* bcd_in1=00101000 bcd_in2=10000011 cout=1 sum=00010001
* bcd_in1=00101000 bcd_in2=10000100 cout=1 sum=00010010
* bcd_in1=00101000 bcd_in2=10000101 cout=1 sum=00010011
* bcd_in1=00101000 bcd_in2=10000110 cout=1 sum=00010100
* bcd_in1=00101000 bcd_in2=10000111 cout=1 sum=00010101
* bcd_in1=00101000 bcd_in2=10001000 cout=1 sum=00010110
* bcd_in1=00101000 bcd_in2=10001001 cout=1 sum=00010111
* bcd_in1=00101000 bcd_in2=10010000 cout=1 sum=00011000
* bcd_in1=00101000 bcd_in2=10010001 cout=1 sum=00011001
* bcd_in1=00101000 bcd_in2=10010010 cout=1 sum=00100000
* bcd_in1=00101000 bcd_in2=10010011 cout=1 sum=00100001
* bcd_in1=00101000 bcd_in2=10010100 cout=1 sum=00100010
* bcd_in1=00101000 bcd_in2=10010101 cout=1 sum=00100011
* bcd_in1=00101000 bcd_in2=10010110 cout=1 sum=00100100
* bcd_in1=00101000 bcd_in2=10010111 cout=1 sum=00100101
* bcd_in1=00101000 bcd_in2=10011000 cout=1 sum=00100110
* bcd_in1=00101000 bcd_in2=10011001 cout=1 sum=00100111
* bcd_in1=00101001 bcd_in2=00000000 cout=0 sum=00101001
* bcd_in1=00101001 bcd_in2=00000001 cout=0 sum=00110000
* bcd_in1=00101001 bcd_in2=00000010 cout=0 sum=00110001
* bcd_in1=00101001 bcd_in2=00000011 cout=0 sum=00110010
* bcd_in1=00101001 bcd_in2=00000100 cout=0 sum=00110011
* bcd_in1=00101001 bcd_in2=00000101 cout=0 sum=00110100
* bcd_in1=00101001 bcd_in2=00000110 cout=0 sum=00110101
* bcd_in1=00101001 bcd_in2=00000111 cout=0 sum=00110110
* bcd_in1=00101001 bcd_in2=00001000 cout=0 sum=00110111
* bcd_in1=00101001 bcd_in2=00001001 cout=0 sum=00111000
* bcd_in1=00101001 bcd_in2=00010000 cout=0 sum=00111001
* bcd_in1=00101001 bcd_in2=00010001 cout=0 sum=01000000
* bcd_in1=00101001 bcd_in2=00010010 cout=0 sum=01000001
* bcd_in1=00101001 bcd_in2=00010011 cout=0 sum=01000010
* bcd_in1=00101001 bcd_in2=00010100 cout=0 sum=01000011
* bcd_in1=00101001 bcd_in2=00010101 cout=0 sum=01000100
* bcd_in1=00101001 bcd_in2=00010110 cout=0 sum=01000101
* bcd_in1=00101001 bcd_in2=00010111 cout=0 sum=01000110
* bcd_in1=00101001 bcd_in2=00011000 cout=0 sum=01000111
* bcd_in1=00101001 bcd_in2=00011001 cout=0 sum=01001000
* bcd_in1=00101001 bcd_in2=00100000 cout=0 sum=01001001
* bcd_in1=00101001 bcd_in2=00100001 cout=0 sum=01010000
* bcd_in1=00101001 bcd_in2=00100010 cout=0 sum=01010001
* bcd_in1=00101001 bcd_in2=00100011 cout=0 sum=01010010
* bcd_in1=00101001 bcd_in2=00100100 cout=0 sum=01010011
* bcd_in1=00101001 bcd_in2=00100101 cout=0 sum=01010100
* bcd_in1=00101001 bcd_in2=00100110 cout=0 sum=01010101
* bcd_in1=00101001 bcd_in2=00100111 cout=0 sum=01010110
* bcd_in1=00101001 bcd_in2=00101000 cout=0 sum=01010111
* bcd_in1=00101001 bcd_in2=00101001 cout=0 sum=01011000
* bcd_in1=00101001 bcd_in2=00110000 cout=0 sum=01011001
* bcd_in1=00101001 bcd_in2=00110001 cout=0 sum=01100000
* bcd_in1=00101001 bcd_in2=00110010 cout=0 sum=01100001
* bcd_in1=00101001 bcd_in2=00110011 cout=0 sum=01100010
* bcd_in1=00101001 bcd_in2=00110100 cout=0 sum=01100011
* bcd_in1=00101001 bcd_in2=00110101 cout=0 sum=01100100
* bcd_in1=00101001 bcd_in2=00110110 cout=0 sum=01100101
* bcd_in1=00101001 bcd_in2=00110111 cout=0 sum=01100110
* bcd_in1=00101001 bcd_in2=00111000 cout=0 sum=01100111
* bcd_in1=00101001 bcd_in2=00111001 cout=0 sum=01101000
* bcd_in1=00101001 bcd_in2=01000000 cout=0 sum=01101001
* bcd_in1=00101001 bcd_in2=01000001 cout=0 sum=01110000
* bcd_in1=00101001 bcd_in2=01000010 cout=0 sum=01110001
* bcd_in1=00101001 bcd_in2=01000011 cout=0 sum=01110010
* bcd_in1=00101001 bcd_in2=01000100 cout=0 sum=01110011
* bcd_in1=00101001 bcd_in2=01000101 cout=0 sum=01110100
* bcd_in1=00101001 bcd_in2=01000110 cout=0 sum=01110101
* bcd_in1=00101001 bcd_in2=01000111 cout=0 sum=01110110
* bcd_in1=00101001 bcd_in2=01001000 cout=0 sum=01110111
* bcd_in1=00101001 bcd_in2=01001001 cout=0 sum=01111000
* bcd_in1=00101001 bcd_in2=01010000 cout=0 sum=01111001
* bcd_in1=00101001 bcd_in2=01010001 cout=0 sum=10000000
* bcd_in1=00101001 bcd_in2=01010010 cout=0 sum=10000001
* bcd_in1=00101001 bcd_in2=01010011 cout=0 sum=10000010
* bcd_in1=00101001 bcd_in2=01010100 cout=0 sum=10000011
* bcd_in1=00101001 bcd_in2=01010101 cout=0 sum=10000100
* bcd_in1=00101001 bcd_in2=01010110 cout=0 sum=10000101
* bcd_in1=00101001 bcd_in2=01010111 cout=0 sum=10000110
* bcd_in1=00101001 bcd_in2=01011000 cout=0 sum=10000111
* bcd_in1=00101001 bcd_in2=01011001 cout=0 sum=10001000
* bcd_in1=00101001 bcd_in2=01100000 cout=0 sum=10001001
* bcd_in1=00101001 bcd_in2=01100001 cout=0 sum=10010000
* bcd_in1=00101001 bcd_in2=01100010 cout=0 sum=10010001
* bcd_in1=00101001 bcd_in2=01100011 cout=0 sum=10010010
* bcd_in1=00101001 bcd_in2=01100100 cout=0 sum=10010011
* bcd_in1=00101001 bcd_in2=01100101 cout=0 sum=10010100
* bcd_in1=00101001 bcd_in2=01100110 cout=0 sum=10010101
* bcd_in1=00101001 bcd_in2=01100111 cout=0 sum=10010110
* bcd_in1=00101001 bcd_in2=01101000 cout=0 sum=10010111
* bcd_in1=00101001 bcd_in2=01101001 cout=0 sum=10011000
* bcd_in1=00101001 bcd_in2=01110000 cout=0 sum=10011001
* bcd_in1=00101001 bcd_in2=01110001 cout=1 sum=00000000
* bcd_in1=00101001 bcd_in2=01110010 cout=1 sum=00000001
* bcd_in1=00101001 bcd_in2=01110011 cout=1 sum=00000010
* bcd_in1=00101001 bcd_in2=01110100 cout=1 sum=00000011
* bcd_in1=00101001 bcd_in2=01110101 cout=1 sum=00000100
* bcd_in1=00101001 bcd_in2=01110110 cout=1 sum=00000101
* bcd_in1=00101001 bcd_in2=01110111 cout=1 sum=00000110
* bcd_in1=00101001 bcd_in2=01111000 cout=1 sum=00000111
* bcd_in1=00101001 bcd_in2=01111001 cout=1 sum=00001000
* bcd_in1=00101001 bcd_in2=10000000 cout=1 sum=00001001
* bcd_in1=00101001 bcd_in2=10000001 cout=1 sum=00010000
* bcd_in1=00101001 bcd_in2=10000010 cout=1 sum=00010001
* bcd_in1=00101001 bcd_in2=10000011 cout=1 sum=00010010
* bcd_in1=00101001 bcd_in2=10000100 cout=1 sum=00010011
* bcd_in1=00101001 bcd_in2=10000101 cout=1 sum=00010100
* bcd_in1=00101001 bcd_in2=10000110 cout=1 sum=00010101
* bcd_in1=00101001 bcd_in2=10000111 cout=1 sum=00010110
* bcd_in1=00101001 bcd_in2=10001000 cout=1 sum=00010111
* bcd_in1=00101001 bcd_in2=10001001 cout=1 sum=00011000
* bcd_in1=00101001 bcd_in2=10010000 cout=1 sum=00011001
* bcd_in1=00101001 bcd_in2=10010001 cout=1 sum=00100000
* bcd_in1=00101001 bcd_in2=10010010 cout=1 sum=00100001
* bcd_in1=00101001 bcd_in2=10010011 cout=1 sum=00100010
* bcd_in1=00101001 bcd_in2=10010100 cout=1 sum=00100011
* bcd_in1=00101001 bcd_in2=10010101 cout=1 sum=00100100
* bcd_in1=00101001 bcd_in2=10010110 cout=1 sum=00100101
* bcd_in1=00101001 bcd_in2=10010111 cout=1 sum=00100110
* bcd_in1=00101001 bcd_in2=10011000 cout=1 sum=00100111
* bcd_in1=00101001 bcd_in2=10011001 cout=1 sum=00101000
* bcd_in1=00110000 bcd_in2=00000000 cout=0 sum=00110000
* bcd_in1=00110000 bcd_in2=00000001 cout=0 sum=00110001
* bcd_in1=00110000 bcd_in2=00000010 cout=0 sum=00110010
* bcd_in1=00110000 bcd_in2=00000011 cout=0 sum=00110011
* bcd_in1=00110000 bcd_in2=00000100 cout=0 sum=00110100
* bcd_in1=00110000 bcd_in2=00000101 cout=0 sum=00110101
* bcd_in1=00110000 bcd_in2=00000110 cout=0 sum=00110110
* bcd_in1=00110000 bcd_in2=00000111 cout=0 sum=00110111
* bcd_in1=00110000 bcd_in2=00001000 cout=0 sum=00111000
* bcd_in1=00110000 bcd_in2=00001001 cout=0 sum=00111001
* bcd_in1=00110000 bcd_in2=00010000 cout=0 sum=01000000
* bcd_in1=00110000 bcd_in2=00010001 cout=0 sum=01000001
* bcd_in1=00110000 bcd_in2=00010010 cout=0 sum=01000010
* bcd_in1=00110000 bcd_in2=00010011 cout=0 sum=01000011
* bcd_in1=00110000 bcd_in2=00010100 cout=0 sum=01000100
* bcd_in1=00110000 bcd_in2=00010101 cout=0 sum=01000101
* bcd_in1=00110000 bcd_in2=00010110 cout=0 sum=01000110
* bcd_in1=00110000 bcd_in2=00010111 cout=0 sum=01000111
* bcd_in1=00110000 bcd_in2=00011000 cout=0 sum=01001000
* bcd_in1=00110000 bcd_in2=00011001 cout=0 sum=01001001
* bcd_in1=00110000 bcd_in2=00100000 cout=0 sum=01010000
* bcd_in1=00110000 bcd_in2=00100001 cout=0 sum=01010001
* bcd_in1=00110000 bcd_in2=00100010 cout=0 sum=01010010
* bcd_in1=00110000 bcd_in2=00100011 cout=0 sum=01010011
* bcd_in1=00110000 bcd_in2=00100100 cout=0 sum=01010100
* bcd_in1=00110000 bcd_in2=00100101 cout=0 sum=01010101
* bcd_in1=00110000 bcd_in2=00100110 cout=0 sum=01010110
* bcd_in1=00110000 bcd_in2=00100111 cout=0 sum=01010111
* bcd_in1=00110000 bcd_in2=00101000 cout=0 sum=01011000
* bcd_in1=00110000 bcd_in2=00101001 cout=0 sum=01011001
* bcd_in1=00110000 bcd_in2=00110000 cout=0 sum=01100000
* bcd_in1=00110000 bcd_in2=00110001 cout=0 sum=01100001
* bcd_in1=00110000 bcd_in2=00110010 cout=0 sum=01100010
* bcd_in1=00110000 bcd_in2=00110011 cout=0 sum=01100011
* bcd_in1=00110000 bcd_in2=00110100 cout=0 sum=01100100
* bcd_in1=00110000 bcd_in2=00110101 cout=0 sum=01100101
* bcd_in1=00110000 bcd_in2=00110110 cout=0 sum=01100110
* bcd_in1=00110000 bcd_in2=00110111 cout=0 sum=01100111
* bcd_in1=00110000 bcd_in2=00111000 cout=0 sum=01101000
* bcd_in1=00110000 bcd_in2=00111001 cout=0 sum=01101001
* bcd_in1=00110000 bcd_in2=01000000 cout=0 sum=01110000
* bcd_in1=00110000 bcd_in2=01000001 cout=0 sum=01110001
* bcd_in1=00110000 bcd_in2=01000010 cout=0 sum=01110010
* bcd_in1=00110000 bcd_in2=01000011 cout=0 sum=01110011
* bcd_in1=00110000 bcd_in2=01000100 cout=0 sum=01110100
* bcd_in1=00110000 bcd_in2=01000101 cout=0 sum=01110101
* bcd_in1=00110000 bcd_in2=01000110 cout=0 sum=01110110
* bcd_in1=00110000 bcd_in2=01000111 cout=0 sum=01110111
* bcd_in1=00110000 bcd_in2=01001000 cout=0 sum=01111000
* bcd_in1=00110000 bcd_in2=01001001 cout=0 sum=01111001
* bcd_in1=00110000 bcd_in2=01010000 cout=0 sum=10000000
* bcd_in1=00110000 bcd_in2=01010001 cout=0 sum=10000001
* bcd_in1=00110000 bcd_in2=01010010 cout=0 sum=10000010
* bcd_in1=00110000 bcd_in2=01010011 cout=0 sum=10000011
* bcd_in1=00110000 bcd_in2=01010100 cout=0 sum=10000100
* bcd_in1=00110000 bcd_in2=01010101 cout=0 sum=10000101
* bcd_in1=00110000 bcd_in2=01010110 cout=0 sum=10000110
* bcd_in1=00110000 bcd_in2=01010111 cout=0 sum=10000111
* bcd_in1=00110000 bcd_in2=01011000 cout=0 sum=10001000
* bcd_in1=00110000 bcd_in2=01011001 cout=0 sum=10001001
* bcd_in1=00110000 bcd_in2=01100000 cout=0 sum=10010000
* bcd_in1=00110000 bcd_in2=01100001 cout=0 sum=10010001
* bcd_in1=00110000 bcd_in2=01100010 cout=0 sum=10010010
* bcd_in1=00110000 bcd_in2=01100011 cout=0 sum=10010011
* bcd_in1=00110000 bcd_in2=01100100 cout=0 sum=10010100
* bcd_in1=00110000 bcd_in2=01100101 cout=0 sum=10010101
* bcd_in1=00110000 bcd_in2=01100110 cout=0 sum=10010110
* bcd_in1=00110000 bcd_in2=01100111 cout=0 sum=10010111
* bcd_in1=00110000 bcd_in2=01101000 cout=0 sum=10011000
* bcd_in1=00110000 bcd_in2=01101001 cout=0 sum=10011001
* bcd_in1=00110000 bcd_in2=01110000 cout=1 sum=00000000
* bcd_in1=00110000 bcd_in2=01110001 cout=1 sum=00000001
* bcd_in1=00110000 bcd_in2=01110010 cout=1 sum=00000010
* bcd_in1=00110000 bcd_in2=01110011 cout=1 sum=00000011
* bcd_in1=00110000 bcd_in2=01110100 cout=1 sum=00000100
* bcd_in1=00110000 bcd_in2=01110101 cout=1 sum=00000101
* bcd_in1=00110000 bcd_in2=01110110 cout=1 sum=00000110
* bcd_in1=00110000 bcd_in2=01110111 cout=1 sum=00000111
* bcd_in1=00110000 bcd_in2=01111000 cout=1 sum=00001000
* bcd_in1=00110000 bcd_in2=01111001 cout=1 sum=00001001
* bcd_in1=00110000 bcd_in2=10000000 cout=1 sum=00010000
* bcd_in1=00110000 bcd_in2=10000001 cout=1 sum=00010001
* bcd_in1=00110000 bcd_in2=10000010 cout=1 sum=00010010
* bcd_in1=00110000 bcd_in2=10000011 cout=1 sum=00010011
* bcd_in1=00110000 bcd_in2=10000100 cout=1 sum=00010100
* bcd_in1=00110000 bcd_in2=10000101 cout=1 sum=00010101
* bcd_in1=00110000 bcd_in2=10000110 cout=1 sum=00010110
* bcd_in1=00110000 bcd_in2=10000111 cout=1 sum=00010111
* bcd_in1=00110000 bcd_in2=10001000 cout=1 sum=00011000
* bcd_in1=00110000 bcd_in2=10001001 cout=1 sum=00011001
* bcd_in1=00110000 bcd_in2=10010000 cout=1 sum=00100000
* bcd_in1=00110000 bcd_in2=10010001 cout=1 sum=00100001
* bcd_in1=00110000 bcd_in2=10010010 cout=1 sum=00100010
* bcd_in1=00110000 bcd_in2=10010011 cout=1 sum=00100011
* bcd_in1=00110000 bcd_in2=10010100 cout=1 sum=00100100
* bcd_in1=00110000 bcd_in2=10010101 cout=1 sum=00100101
* bcd_in1=00110000 bcd_in2=10010110 cout=1 sum=00100110
* bcd_in1=00110000 bcd_in2=10010111 cout=1 sum=00100111
* bcd_in1=00110000 bcd_in2=10011000 cout=1 sum=00101000
* bcd_in1=00110000 bcd_in2=10011001 cout=1 sum=00101001
* bcd_in1=00110001 bcd_in2=00000000 cout=0 sum=00110001
* bcd_in1=00110001 bcd_in2=00000001 cout=0 sum=00110010
* bcd_in1=00110001 bcd_in2=00000010 cout=0 sum=00110011
* bcd_in1=00110001 bcd_in2=00000011 cout=0 sum=00110100
* bcd_in1=00110001 bcd_in2=00000100 cout=0 sum=00110101
* bcd_in1=00110001 bcd_in2=00000101 cout=0 sum=00110110
* bcd_in1=00110001 bcd_in2=00000110 cout=0 sum=00110111
* bcd_in1=00110001 bcd_in2=00000111 cout=0 sum=00111000
* bcd_in1=00110001 bcd_in2=00001000 cout=0 sum=00111001
* bcd_in1=00110001 bcd_in2=00001001 cout=0 sum=01000000
* bcd_in1=00110001 bcd_in2=00010000 cout=0 sum=01000001
* bcd_in1=00110001 bcd_in2=00010001 cout=0 sum=01000010
* bcd_in1=00110001 bcd_in2=00010010 cout=0 sum=01000011
* bcd_in1=00110001 bcd_in2=00010011 cout=0 sum=01000100
* bcd_in1=00110001 bcd_in2=00010100 cout=0 sum=01000101
* bcd_in1=00110001 bcd_in2=00010101 cout=0 sum=01000110
* bcd_in1=00110001 bcd_in2=00010110 cout=0 sum=01000111
* bcd_in1=00110001 bcd_in2=00010111 cout=0 sum=01001000
* bcd_in1=00110001 bcd_in2=00011000 cout=0 sum=01001001
* bcd_in1=00110001 bcd_in2=00011001 cout=0 sum=01010000
* bcd_in1=00110001 bcd_in2=00100000 cout=0 sum=01010001
* bcd_in1=00110001 bcd_in2=00100001 cout=0 sum=01010010
* bcd_in1=00110001 bcd_in2=00100010 cout=0 sum=01010011
* bcd_in1=00110001 bcd_in2=00100011 cout=0 sum=01010100
* bcd_in1=00110001 bcd_in2=00100100 cout=0 sum=01010101
* bcd_in1=00110001 bcd_in2=00100101 cout=0 sum=01010110
* bcd_in1=00110001 bcd_in2=00100110 cout=0 sum=01010111
* bcd_in1=00110001 bcd_in2=00100111 cout=0 sum=01011000
* bcd_in1=00110001 bcd_in2=00101000 cout=0 sum=01011001
* bcd_in1=00110001 bcd_in2=00101001 cout=0 sum=01100000
* bcd_in1=00110001 bcd_in2=00110000 cout=0 sum=01100001
* bcd_in1=00110001 bcd_in2=00110001 cout=0 sum=01100010
* bcd_in1=00110001 bcd_in2=00110010 cout=0 sum=01100011
* bcd_in1=00110001 bcd_in2=00110011 cout=0 sum=01100100
* bcd_in1=00110001 bcd_in2=00110100 cout=0 sum=01100101
* bcd_in1=00110001 bcd_in2=00110101 cout=0 sum=01100110
* bcd_in1=00110001 bcd_in2=00110110 cout=0 sum=01100111
* bcd_in1=00110001 bcd_in2=00110111 cout=0 sum=01101000
* bcd_in1=00110001 bcd_in2=00111000 cout=0 sum=01101001
* bcd_in1=00110001 bcd_in2=00111001 cout=0 sum=01110000
* bcd_in1=00110001 bcd_in2=01000000 cout=0 sum=01110001
* bcd_in1=00110001 bcd_in2=01000001 cout=0 sum=01110010
* bcd_in1=00110001 bcd_in2=01000010 cout=0 sum=01110011
* bcd_in1=00110001 bcd_in2=01000011 cout=0 sum=01110100
* bcd_in1=00110001 bcd_in2=01000100 cout=0 sum=01110101
* bcd_in1=00110001 bcd_in2=01000101 cout=0 sum=01110110
* bcd_in1=00110001 bcd_in2=01000110 cout=0 sum=01110111
* bcd_in1=00110001 bcd_in2=01000111 cout=0 sum=01111000
* bcd_in1=00110001 bcd_in2=01001000 cout=0 sum=01111001
* bcd_in1=00110001 bcd_in2=01001001 cout=0 sum=10000000
* bcd_in1=00110001 bcd_in2=01010000 cout=0 sum=10000001
* bcd_in1=00110001 bcd_in2=01010001 cout=0 sum=10000010
* bcd_in1=00110001 bcd_in2=01010010 cout=0 sum=10000011
* bcd_in1=00110001 bcd_in2=01010011 cout=0 sum=10000100
* bcd_in1=00110001 bcd_in2=01010100 cout=0 sum=10000101
* bcd_in1=00110001 bcd_in2=01010101 cout=0 sum=10000110
* bcd_in1=00110001 bcd_in2=01010110 cout=0 sum=10000111
* bcd_in1=00110001 bcd_in2=01010111 cout=0 sum=10001000
* bcd_in1=00110001 bcd_in2=01011000 cout=0 sum=10001001
* bcd_in1=00110001 bcd_in2=01011001 cout=0 sum=10010000
* bcd_in1=00110001 bcd_in2=01100000 cout=0 sum=10010001
* bcd_in1=00110001 bcd_in2=01100001 cout=0 sum=10010010
* bcd_in1=00110001 bcd_in2=01100010 cout=0 sum=10010011
* bcd_in1=00110001 bcd_in2=01100011 cout=0 sum=10010100
* bcd_in1=00110001 bcd_in2=01100100 cout=0 sum=10010101
* bcd_in1=00110001 bcd_in2=01100101 cout=0 sum=10010110
* bcd_in1=00110001 bcd_in2=01100110 cout=0 sum=10010111
* bcd_in1=00110001 bcd_in2=01100111 cout=0 sum=10011000
* bcd_in1=00110001 bcd_in2=01101000 cout=0 sum=10011001
* bcd_in1=00110001 bcd_in2=01101001 cout=1 sum=00000000
* bcd_in1=00110001 bcd_in2=01110000 cout=1 sum=00000001
* bcd_in1=00110001 bcd_in2=01110001 cout=1 sum=00000010
* bcd_in1=00110001 bcd_in2=01110010 cout=1 sum=00000011
* bcd_in1=00110001 bcd_in2=01110011 cout=1 sum=00000100
* bcd_in1=00110001 bcd_in2=01110100 cout=1 sum=00000101
* bcd_in1=00110001 bcd_in2=01110101 cout=1 sum=00000110
* bcd_in1=00110001 bcd_in2=01110110 cout=1 sum=00000111
* bcd_in1=00110001 bcd_in2=01110111 cout=1 sum=00001000
* bcd_in1=00110001 bcd_in2=01111000 cout=1 sum=00001001
* bcd_in1=00110001 bcd_in2=01111001 cout=1 sum=00010000
* bcd_in1=00110001 bcd_in2=10000000 cout=1 sum=00010001
* bcd_in1=00110001 bcd_in2=10000001 cout=1 sum=00010010
* bcd_in1=00110001 bcd_in2=10000010 cout=1 sum=00010011
* bcd_in1=00110001 bcd_in2=10000011 cout=1 sum=00010100
* bcd_in1=00110001 bcd_in2=10000100 cout=1 sum=00010101
* bcd_in1=00110001 bcd_in2=10000101 cout=1 sum=00010110
* bcd_in1=00110001 bcd_in2=10000110 cout=1 sum=00010111
* bcd_in1=00110001 bcd_in2=10000111 cout=1 sum=00011000
* bcd_in1=00110001 bcd_in2=10001000 cout=1 sum=00011001
* bcd_in1=00110001 bcd_in2=10001001 cout=1 sum=00100000
* bcd_in1=00110001 bcd_in2=10010000 cout=1 sum=00100001
* bcd_in1=00110001 bcd_in2=10010001 cout=1 sum=00100010
* bcd_in1=00110001 bcd_in2=10010010 cout=1 sum=00100011
* bcd_in1=00110001 bcd_in2=10010011 cout=1 sum=00100100
* bcd_in1=00110001 bcd_in2=10010100 cout=1 sum=00100101
* bcd_in1=00110001 bcd_in2=10010101 cout=1 sum=00100110
* bcd_in1=00110001 bcd_in2=10010110 cout=1 sum=00100111
* bcd_in1=00110001 bcd_in2=10010111 cout=1 sum=00101000
* bcd_in1=00110001 bcd_in2=10011000 cout=1 sum=00101001
* bcd_in1=00110001 bcd_in2=10011001 cout=1 sum=00110000
* bcd_in1=00110010 bcd_in2=00000000 cout=0 sum=00110010
* bcd_in1=00110010 bcd_in2=00000001 cout=0 sum=00110011
* bcd_in1=00110010 bcd_in2=00000010 cout=0 sum=00110100
* bcd_in1=00110010 bcd_in2=00000011 cout=0 sum=00110101
* bcd_in1=00110010 bcd_in2=00000100 cout=0 sum=00110110
* bcd_in1=00110010 bcd_in2=00000101 cout=0 sum=00110111
* bcd_in1=00110010 bcd_in2=00000110 cout=0 sum=00111000
* bcd_in1=00110010 bcd_in2=00000111 cout=0 sum=00111001
* bcd_in1=00110010 bcd_in2=00001000 cout=0 sum=01000000
* bcd_in1=00110010 bcd_in2=00001001 cout=0 sum=01000001
* bcd_in1=00110010 bcd_in2=00010000 cout=0 sum=01000010
* bcd_in1=00110010 bcd_in2=00010001 cout=0 sum=01000011
* bcd_in1=00110010 bcd_in2=00010010 cout=0 sum=01000100
* bcd_in1=00110010 bcd_in2=00010011 cout=0 sum=01000101
* bcd_in1=00110010 bcd_in2=00010100 cout=0 sum=01000110
* bcd_in1=00110010 bcd_in2=00010101 cout=0 sum=01000111
* bcd_in1=00110010 bcd_in2=00010110 cout=0 sum=01001000
* bcd_in1=00110010 bcd_in2=00010111 cout=0 sum=01001001
* bcd_in1=00110010 bcd_in2=00011000 cout=0 sum=01010000
* bcd_in1=00110010 bcd_in2=00011001 cout=0 sum=01010001
* bcd_in1=00110010 bcd_in2=00100000 cout=0 sum=01010010
* bcd_in1=00110010 bcd_in2=00100001 cout=0 sum=01010011
* bcd_in1=00110010 bcd_in2=00100010 cout=0 sum=01010100
* bcd_in1=00110010 bcd_in2=00100011 cout=0 sum=01010101
* bcd_in1=00110010 bcd_in2=00100100 cout=0 sum=01010110
* bcd_in1=00110010 bcd_in2=00100101 cout=0 sum=01010111
* bcd_in1=00110010 bcd_in2=00100110 cout=0 sum=01011000
* bcd_in1=00110010 bcd_in2=00100111 cout=0 sum=01011001
* bcd_in1=00110010 bcd_in2=00101000 cout=0 sum=01100000
* bcd_in1=00110010 bcd_in2=00101001 cout=0 sum=01100001
* bcd_in1=00110010 bcd_in2=00110000 cout=0 sum=01100010
* bcd_in1=00110010 bcd_in2=00110001 cout=0 sum=01100011
* bcd_in1=00110010 bcd_in2=00110010 cout=0 sum=01100100
* bcd_in1=00110010 bcd_in2=00110011 cout=0 sum=01100101
* bcd_in1=00110010 bcd_in2=00110100 cout=0 sum=01100110
* bcd_in1=00110010 bcd_in2=00110101 cout=0 sum=01100111
* bcd_in1=00110010 bcd_in2=00110110 cout=0 sum=01101000
* bcd_in1=00110010 bcd_in2=00110111 cout=0 sum=01101001
* bcd_in1=00110010 bcd_in2=00111000 cout=0 sum=01110000
* bcd_in1=00110010 bcd_in2=00111001 cout=0 sum=01110001
* bcd_in1=00110010 bcd_in2=01000000 cout=0 sum=01110010
* bcd_in1=00110010 bcd_in2=01000001 cout=0 sum=01110011
* bcd_in1=00110010 bcd_in2=01000010 cout=0 sum=01110100
* bcd_in1=00110010 bcd_in2=01000011 cout=0 sum=01110101
* bcd_in1=00110010 bcd_in2=01000100 cout=0 sum=01110110
* bcd_in1=00110010 bcd_in2=01000101 cout=0 sum=01110111
* bcd_in1=00110010 bcd_in2=01000110 cout=0 sum=01111000
* bcd_in1=00110010 bcd_in2=01000111 cout=0 sum=01111001
* bcd_in1=00110010 bcd_in2=01001000 cout=0 sum=10000000
* bcd_in1=00110010 bcd_in2=01001001 cout=0 sum=10000001
* bcd_in1=00110010 bcd_in2=01010000 cout=0 sum=10000010
* bcd_in1=00110010 bcd_in2=01010001 cout=0 sum=10000011
* bcd_in1=00110010 bcd_in2=01010010 cout=0 sum=10000100
* bcd_in1=00110010 bcd_in2=01010011 cout=0 sum=10000101
* bcd_in1=00110010 bcd_in2=01010100 cout=0 sum=10000110
* bcd_in1=00110010 bcd_in2=01010101 cout=0 sum=10000111
* bcd_in1=00110010 bcd_in2=01010110 cout=0 sum=10001000
* bcd_in1=00110010 bcd_in2=01010111 cout=0 sum=10001001
* bcd_in1=00110010 bcd_in2=01011000 cout=0 sum=10010000
* bcd_in1=00110010 bcd_in2=01011001 cout=0 sum=10010001
* bcd_in1=00110010 bcd_in2=01100000 cout=0 sum=10010010
* bcd_in1=00110010 bcd_in2=01100001 cout=0 sum=10010011
* bcd_in1=00110010 bcd_in2=01100010 cout=0 sum=10010100
* bcd_in1=00110010 bcd_in2=01100011 cout=0 sum=10010101
* bcd_in1=00110010 bcd_in2=01100100 cout=0 sum=10010110
* bcd_in1=00110010 bcd_in2=01100101 cout=0 sum=10010111
* bcd_in1=00110010 bcd_in2=01100110 cout=0 sum=10011000
* bcd_in1=00110010 bcd_in2=01100111 cout=0 sum=10011001
* bcd_in1=00110010 bcd_in2=01101000 cout=1 sum=00000000
* bcd_in1=00110010 bcd_in2=01101001 cout=1 sum=00000001
* bcd_in1=00110010 bcd_in2=01110000 cout=1 sum=00000010
* bcd_in1=00110010 bcd_in2=01110001 cout=1 sum=00000011
* bcd_in1=00110010 bcd_in2=01110010 cout=1 sum=00000100
* bcd_in1=00110010 bcd_in2=01110011 cout=1 sum=00000101
* bcd_in1=00110010 bcd_in2=01110100 cout=1 sum=00000110
* bcd_in1=00110010 bcd_in2=01110101 cout=1 sum=00000111
* bcd_in1=00110010 bcd_in2=01110110 cout=1 sum=00001000
* bcd_in1=00110010 bcd_in2=01110111 cout=1 sum=00001001
* bcd_in1=00110010 bcd_in2=01111000 cout=1 sum=00010000
* bcd_in1=00110010 bcd_in2=01111001 cout=1 sum=00010001
* bcd_in1=00110010 bcd_in2=10000000 cout=1 sum=00010010
* bcd_in1=00110010 bcd_in2=10000001 cout=1 sum=00010011
* bcd_in1=00110010 bcd_in2=10000010 cout=1 sum=00010100
* bcd_in1=00110010 bcd_in2=10000011 cout=1 sum=00010101
* bcd_in1=00110010 bcd_in2=10000100 cout=1 sum=00010110
* bcd_in1=00110010 bcd_in2=10000101 cout=1 sum=00010111
* bcd_in1=00110010 bcd_in2=10000110 cout=1 sum=00011000
* bcd_in1=00110010 bcd_in2=10000111 cout=1 sum=00011001
* bcd_in1=00110010 bcd_in2=10001000 cout=1 sum=00100000
* bcd_in1=00110010 bcd_in2=10001001 cout=1 sum=00100001
* bcd_in1=00110010 bcd_in2=10010000 cout=1 sum=00100010
* bcd_in1=00110010 bcd_in2=10010001 cout=1 sum=00100011
* bcd_in1=00110010 bcd_in2=10010010 cout=1 sum=00100100
* bcd_in1=00110010 bcd_in2=10010011 cout=1 sum=00100101
* bcd_in1=00110010 bcd_in2=10010100 cout=1 sum=00100110
* bcd_in1=00110010 bcd_in2=10010101 cout=1 sum=00100111
* bcd_in1=00110010 bcd_in2=10010110 cout=1 sum=00101000
* bcd_in1=00110010 bcd_in2=10010111 cout=1 sum=00101001
* bcd_in1=00110010 bcd_in2=10011000 cout=1 sum=00110000
* bcd_in1=00110010 bcd_in2=10011001 cout=1 sum=00110001
* bcd_in1=00110011 bcd_in2=00000000 cout=0 sum=00110011
* bcd_in1=00110011 bcd_in2=00000001 cout=0 sum=00110100
* bcd_in1=00110011 bcd_in2=00000010 cout=0 sum=00110101
* bcd_in1=00110011 bcd_in2=00000011 cout=0 sum=00110110
* bcd_in1=00110011 bcd_in2=00000100 cout=0 sum=00110111
* bcd_in1=00110011 bcd_in2=00000101 cout=0 sum=00111000
* bcd_in1=00110011 bcd_in2=00000110 cout=0 sum=00111001
* bcd_in1=00110011 bcd_in2=00000111 cout=0 sum=01000000
* bcd_in1=00110011 bcd_in2=00001000 cout=0 sum=01000001
* bcd_in1=00110011 bcd_in2=00001001 cout=0 sum=01000010
* bcd_in1=00110011 bcd_in2=00010000 cout=0 sum=01000011
* bcd_in1=00110011 bcd_in2=00010001 cout=0 sum=01000100
* bcd_in1=00110011 bcd_in2=00010010 cout=0 sum=01000101
* bcd_in1=00110011 bcd_in2=00010011 cout=0 sum=01000110
* bcd_in1=00110011 bcd_in2=00010100 cout=0 sum=01000111
* bcd_in1=00110011 bcd_in2=00010101 cout=0 sum=01001000
* bcd_in1=00110011 bcd_in2=00010110 cout=0 sum=01001001
* bcd_in1=00110011 bcd_in2=00010111 cout=0 sum=01010000
* bcd_in1=00110011 bcd_in2=00011000 cout=0 sum=01010001
* bcd_in1=00110011 bcd_in2=00011001 cout=0 sum=01010010
* bcd_in1=00110011 bcd_in2=00100000 cout=0 sum=01010011
* bcd_in1=00110011 bcd_in2=00100001 cout=0 sum=01010100
* bcd_in1=00110011 bcd_in2=00100010 cout=0 sum=01010101
* bcd_in1=00110011 bcd_in2=00100011 cout=0 sum=01010110
* bcd_in1=00110011 bcd_in2=00100100 cout=0 sum=01010111
* bcd_in1=00110011 bcd_in2=00100101 cout=0 sum=01011000
* bcd_in1=00110011 bcd_in2=00100110 cout=0 sum=01011001
* bcd_in1=00110011 bcd_in2=00100111 cout=0 sum=01100000
* bcd_in1=00110011 bcd_in2=00101000 cout=0 sum=01100001
* bcd_in1=00110011 bcd_in2=00101001 cout=0 sum=01100010
* bcd_in1=00110011 bcd_in2=00110000 cout=0 sum=01100011
* bcd_in1=00110011 bcd_in2=00110001 cout=0 sum=01100100
* bcd_in1=00110011 bcd_in2=00110010 cout=0 sum=01100101
* bcd_in1=00110011 bcd_in2=00110011 cout=0 sum=01100110
* bcd_in1=00110011 bcd_in2=00110100 cout=0 sum=01100111
* bcd_in1=00110011 bcd_in2=00110101 cout=0 sum=01101000
* bcd_in1=00110011 bcd_in2=00110110 cout=0 sum=01101001
* bcd_in1=00110011 bcd_in2=00110111 cout=0 sum=01110000
* bcd_in1=00110011 bcd_in2=00111000 cout=0 sum=01110001
* bcd_in1=00110011 bcd_in2=00111001 cout=0 sum=01110010
* bcd_in1=00110011 bcd_in2=01000000 cout=0 sum=01110011
* bcd_in1=00110011 bcd_in2=01000001 cout=0 sum=01110100
* bcd_in1=00110011 bcd_in2=01000010 cout=0 sum=01110101
* bcd_in1=00110011 bcd_in2=01000011 cout=0 sum=01110110
* bcd_in1=00110011 bcd_in2=01000100 cout=0 sum=01110111
* bcd_in1=00110011 bcd_in2=01000101 cout=0 sum=01111000
* bcd_in1=00110011 bcd_in2=01000110 cout=0 sum=01111001
* bcd_in1=00110011 bcd_in2=01000111 cout=0 sum=10000000
* bcd_in1=00110011 bcd_in2=01001000 cout=0 sum=10000001
* bcd_in1=00110011 bcd_in2=01001001 cout=0 sum=10000010
* bcd_in1=00110011 bcd_in2=01010000 cout=0 sum=10000011
* bcd_in1=00110011 bcd_in2=01010001 cout=0 sum=10000100
* bcd_in1=00110011 bcd_in2=01010010 cout=0 sum=10000101
* bcd_in1=00110011 bcd_in2=01010011 cout=0 sum=10000110
* bcd_in1=00110011 bcd_in2=01010100 cout=0 sum=10000111
* bcd_in1=00110011 bcd_in2=01010101 cout=0 sum=10001000
* bcd_in1=00110011 bcd_in2=01010110 cout=0 sum=10001001
* bcd_in1=00110011 bcd_in2=01010111 cout=0 sum=10010000
* bcd_in1=00110011 bcd_in2=01011000 cout=0 sum=10010001
* bcd_in1=00110011 bcd_in2=01011001 cout=0 sum=10010010
* bcd_in1=00110011 bcd_in2=01100000 cout=0 sum=10010011
* bcd_in1=00110011 bcd_in2=01100001 cout=0 sum=10010100
* bcd_in1=00110011 bcd_in2=01100010 cout=0 sum=10010101
* bcd_in1=00110011 bcd_in2=01100011 cout=0 sum=10010110
* bcd_in1=00110011 bcd_in2=01100100 cout=0 sum=10010111
* bcd_in1=00110011 bcd_in2=01100101 cout=0 sum=10011000
* bcd_in1=00110011 bcd_in2=01100110 cout=0 sum=10011001
* bcd_in1=00110011 bcd_in2=01100111 cout=1 sum=00000000
* bcd_in1=00110011 bcd_in2=01101000 cout=1 sum=00000001
* bcd_in1=00110011 bcd_in2=01101001 cout=1 sum=00000010
* bcd_in1=00110011 bcd_in2=01110000 cout=1 sum=00000011
* bcd_in1=00110011 bcd_in2=01110001 cout=1 sum=00000100
* bcd_in1=00110011 bcd_in2=01110010 cout=1 sum=00000101
* bcd_in1=00110011 bcd_in2=01110011 cout=1 sum=00000110
* bcd_in1=00110011 bcd_in2=01110100 cout=1 sum=00000111
* bcd_in1=00110011 bcd_in2=01110101 cout=1 sum=00001000
* bcd_in1=00110011 bcd_in2=01110110 cout=1 sum=00001001
* bcd_in1=00110011 bcd_in2=01110111 cout=1 sum=00010000
* bcd_in1=00110011 bcd_in2=01111000 cout=1 sum=00010001
* bcd_in1=00110011 bcd_in2=01111001 cout=1 sum=00010010
* bcd_in1=00110011 bcd_in2=10000000 cout=1 sum=00010011
* bcd_in1=00110011 bcd_in2=10000001 cout=1 sum=00010100
* bcd_in1=00110011 bcd_in2=10000010 cout=1 sum=00010101
* bcd_in1=00110011 bcd_in2=10000011 cout=1 sum=00010110
* bcd_in1=00110011 bcd_in2=10000100 cout=1 sum=00010111
* bcd_in1=00110011 bcd_in2=10000101 cout=1 sum=00011000
* bcd_in1=00110011 bcd_in2=10000110 cout=1 sum=00011001
* bcd_in1=00110011 bcd_in2=10000111 cout=1 sum=00100000
* bcd_in1=00110011 bcd_in2=10001000 cout=1 sum=00100001
* bcd_in1=00110011 bcd_in2=10001001 cout=1 sum=00100010
* bcd_in1=00110011 bcd_in2=10010000 cout=1 sum=00100011
* bcd_in1=00110011 bcd_in2=10010001 cout=1 sum=00100100
* bcd_in1=00110011 bcd_in2=10010010 cout=1 sum=00100101
* bcd_in1=00110011 bcd_in2=10010011 cout=1 sum=00100110
* bcd_in1=00110011 bcd_in2=10010100 cout=1 sum=00100111
* bcd_in1=00110011 bcd_in2=10010101 cout=1 sum=00101000
* bcd_in1=00110011 bcd_in2=10010110 cout=1 sum=00101001
* bcd_in1=00110011 bcd_in2=10010111 cout=1 sum=00110000
* bcd_in1=00110011 bcd_in2=10011000 cout=1 sum=00110001
* bcd_in1=00110011 bcd_in2=10011001 cout=1 sum=00110010
* bcd_in1=00110100 bcd_in2=00000000 cout=0 sum=00110100
* bcd_in1=00110100 bcd_in2=00000001 cout=0 sum=00110101
* bcd_in1=00110100 bcd_in2=00000010 cout=0 sum=00110110
* bcd_in1=00110100 bcd_in2=00000011 cout=0 sum=00110111
* bcd_in1=00110100 bcd_in2=00000100 cout=0 sum=00111000
* bcd_in1=00110100 bcd_in2=00000101 cout=0 sum=00111001
* bcd_in1=00110100 bcd_in2=00000110 cout=0 sum=01000000
* bcd_in1=00110100 bcd_in2=00000111 cout=0 sum=01000001
* bcd_in1=00110100 bcd_in2=00001000 cout=0 sum=01000010
* bcd_in1=00110100 bcd_in2=00001001 cout=0 sum=01000011
* bcd_in1=00110100 bcd_in2=00010000 cout=0 sum=01000100
* bcd_in1=00110100 bcd_in2=00010001 cout=0 sum=01000101
* bcd_in1=00110100 bcd_in2=00010010 cout=0 sum=01000110
* bcd_in1=00110100 bcd_in2=00010011 cout=0 sum=01000111
* bcd_in1=00110100 bcd_in2=00010100 cout=0 sum=01001000
* bcd_in1=00110100 bcd_in2=00010101 cout=0 sum=01001001
* bcd_in1=00110100 bcd_in2=00010110 cout=0 sum=01010000
* bcd_in1=00110100 bcd_in2=00010111 cout=0 sum=01010001
* bcd_in1=00110100 bcd_in2=00011000 cout=0 sum=01010010
* bcd_in1=00110100 bcd_in2=00011001 cout=0 sum=01010011
* bcd_in1=00110100 bcd_in2=00100000 cout=0 sum=01010100
* bcd_in1=00110100 bcd_in2=00100001 cout=0 sum=01010101
* bcd_in1=00110100 bcd_in2=00100010 cout=0 sum=01010110
* bcd_in1=00110100 bcd_in2=00100011 cout=0 sum=01010111
* bcd_in1=00110100 bcd_in2=00100100 cout=0 sum=01011000
* bcd_in1=00110100 bcd_in2=00100101 cout=0 sum=01011001
* bcd_in1=00110100 bcd_in2=00100110 cout=0 sum=01100000
* bcd_in1=00110100 bcd_in2=00100111 cout=0 sum=01100001
* bcd_in1=00110100 bcd_in2=00101000 cout=0 sum=01100010
* bcd_in1=00110100 bcd_in2=00101001 cout=0 sum=01100011
* bcd_in1=00110100 bcd_in2=00110000 cout=0 sum=01100100
* bcd_in1=00110100 bcd_in2=00110001 cout=0 sum=01100101
* bcd_in1=00110100 bcd_in2=00110010 cout=0 sum=01100110
* bcd_in1=00110100 bcd_in2=00110011 cout=0 sum=01100111
* bcd_in1=00110100 bcd_in2=00110100 cout=0 sum=01101000
* bcd_in1=00110100 bcd_in2=00110101 cout=0 sum=01101001
* bcd_in1=00110100 bcd_in2=00110110 cout=0 sum=01110000
* bcd_in1=00110100 bcd_in2=00110111 cout=0 sum=01110001
* bcd_in1=00110100 bcd_in2=00111000 cout=0 sum=01110010
* bcd_in1=00110100 bcd_in2=00111001 cout=0 sum=01110011
* bcd_in1=00110100 bcd_in2=01000000 cout=0 sum=01110100
* bcd_in1=00110100 bcd_in2=01000001 cout=0 sum=01110101
* bcd_in1=00110100 bcd_in2=01000010 cout=0 sum=01110110
* bcd_in1=00110100 bcd_in2=01000011 cout=0 sum=01110111
* bcd_in1=00110100 bcd_in2=01000100 cout=0 sum=01111000
* bcd_in1=00110100 bcd_in2=01000101 cout=0 sum=01111001
* bcd_in1=00110100 bcd_in2=01000110 cout=0 sum=10000000
* bcd_in1=00110100 bcd_in2=01000111 cout=0 sum=10000001
* bcd_in1=00110100 bcd_in2=01001000 cout=0 sum=10000010
* bcd_in1=00110100 bcd_in2=01001001 cout=0 sum=10000011
* bcd_in1=00110100 bcd_in2=01010000 cout=0 sum=10000100
* bcd_in1=00110100 bcd_in2=01010001 cout=0 sum=10000101
* bcd_in1=00110100 bcd_in2=01010010 cout=0 sum=10000110
* bcd_in1=00110100 bcd_in2=01010011 cout=0 sum=10000111
* bcd_in1=00110100 bcd_in2=01010100 cout=0 sum=10001000
* bcd_in1=00110100 bcd_in2=01010101 cout=0 sum=10001001
* bcd_in1=00110100 bcd_in2=01010110 cout=0 sum=10010000
* bcd_in1=00110100 bcd_in2=01010111 cout=0 sum=10010001
* bcd_in1=00110100 bcd_in2=01011000 cout=0 sum=10010010
* bcd_in1=00110100 bcd_in2=01011001 cout=0 sum=10010011
* bcd_in1=00110100 bcd_in2=01100000 cout=0 sum=10010100
* bcd_in1=00110100 bcd_in2=01100001 cout=0 sum=10010101
* bcd_in1=00110100 bcd_in2=01100010 cout=0 sum=10010110
* bcd_in1=00110100 bcd_in2=01100011 cout=0 sum=10010111
* bcd_in1=00110100 bcd_in2=01100100 cout=0 sum=10011000
* bcd_in1=00110100 bcd_in2=01100101 cout=0 sum=10011001
* bcd_in1=00110100 bcd_in2=01100110 cout=1 sum=00000000
* bcd_in1=00110100 bcd_in2=01100111 cout=1 sum=00000001
* bcd_in1=00110100 bcd_in2=01101000 cout=1 sum=00000010
* bcd_in1=00110100 bcd_in2=01101001 cout=1 sum=00000011
* bcd_in1=00110100 bcd_in2=01110000 cout=1 sum=00000100
* bcd_in1=00110100 bcd_in2=01110001 cout=1 sum=00000101
* bcd_in1=00110100 bcd_in2=01110010 cout=1 sum=00000110
* bcd_in1=00110100 bcd_in2=01110011 cout=1 sum=00000111
* bcd_in1=00110100 bcd_in2=01110100 cout=1 sum=00001000
* bcd_in1=00110100 bcd_in2=01110101 cout=1 sum=00001001
* bcd_in1=00110100 bcd_in2=01110110 cout=1 sum=00010000
* bcd_in1=00110100 bcd_in2=01110111 cout=1 sum=00010001
* bcd_in1=00110100 bcd_in2=01111000 cout=1 sum=00010010
* bcd_in1=00110100 bcd_in2=01111001 cout=1 sum=00010011
* bcd_in1=00110100 bcd_in2=10000000 cout=1 sum=00010100
* bcd_in1=00110100 bcd_in2=10000001 cout=1 sum=00010101
* bcd_in1=00110100 bcd_in2=10000010 cout=1 sum=00010110
* bcd_in1=00110100 bcd_in2=10000011 cout=1 sum=00010111
* bcd_in1=00110100 bcd_in2=10000100 cout=1 sum=00011000
* bcd_in1=00110100 bcd_in2=10000101 cout=1 sum=00011001
* bcd_in1=00110100 bcd_in2=10000110 cout=1 sum=00100000
* bcd_in1=00110100 bcd_in2=10000111 cout=1 sum=00100001
* bcd_in1=00110100 bcd_in2=10001000 cout=1 sum=00100010
* bcd_in1=00110100 bcd_in2=10001001 cout=1 sum=00100011
* bcd_in1=00110100 bcd_in2=10010000 cout=1 sum=00100100
* bcd_in1=00110100 bcd_in2=10010001 cout=1 sum=00100101
* bcd_in1=00110100 bcd_in2=10010010 cout=1 sum=00100110
* bcd_in1=00110100 bcd_in2=10010011 cout=1 sum=00100111
* bcd_in1=00110100 bcd_in2=10010100 cout=1 sum=00101000
* bcd_in1=00110100 bcd_in2=10010101 cout=1 sum=00101001
* bcd_in1=00110100 bcd_in2=10010110 cout=1 sum=00110000
* bcd_in1=00110100 bcd_in2=10010111 cout=1 sum=00110001
* bcd_in1=00110100 bcd_in2=10011000 cout=1 sum=00110010
* bcd_in1=00110100 bcd_in2=10011001 cout=1 sum=00110011
* bcd_in1=00110101 bcd_in2=00000000 cout=0 sum=00110101
* bcd_in1=00110101 bcd_in2=00000001 cout=0 sum=00110110
* bcd_in1=00110101 bcd_in2=00000010 cout=0 sum=00110111
* bcd_in1=00110101 bcd_in2=00000011 cout=0 sum=00111000
* bcd_in1=00110101 bcd_in2=00000100 cout=0 sum=00111001
* bcd_in1=00110101 bcd_in2=00000101 cout=0 sum=01000000
* bcd_in1=00110101 bcd_in2=00000110 cout=0 sum=01000001
* bcd_in1=00110101 bcd_in2=00000111 cout=0 sum=01000010
* bcd_in1=00110101 bcd_in2=00001000 cout=0 sum=01000011
* bcd_in1=00110101 bcd_in2=00001001 cout=0 sum=01000100
* bcd_in1=00110101 bcd_in2=00010000 cout=0 sum=01000101
* bcd_in1=00110101 bcd_in2=00010001 cout=0 sum=01000110
* bcd_in1=00110101 bcd_in2=00010010 cout=0 sum=01000111
* bcd_in1=00110101 bcd_in2=00010011 cout=0 sum=01001000
* bcd_in1=00110101 bcd_in2=00010100 cout=0 sum=01001001
* bcd_in1=00110101 bcd_in2=00010101 cout=0 sum=01010000
* bcd_in1=00110101 bcd_in2=00010110 cout=0 sum=01010001
* bcd_in1=00110101 bcd_in2=00010111 cout=0 sum=01010010
* bcd_in1=00110101 bcd_in2=00011000 cout=0 sum=01010011
* bcd_in1=00110101 bcd_in2=00011001 cout=0 sum=01010100
* bcd_in1=00110101 bcd_in2=00100000 cout=0 sum=01010101
* bcd_in1=00110101 bcd_in2=00100001 cout=0 sum=01010110
* bcd_in1=00110101 bcd_in2=00100010 cout=0 sum=01010111
* bcd_in1=00110101 bcd_in2=00100011 cout=0 sum=01011000
* bcd_in1=00110101 bcd_in2=00100100 cout=0 sum=01011001
* bcd_in1=00110101 bcd_in2=00100101 cout=0 sum=01100000
* bcd_in1=00110101 bcd_in2=00100110 cout=0 sum=01100001
* bcd_in1=00110101 bcd_in2=00100111 cout=0 sum=01100010
* bcd_in1=00110101 bcd_in2=00101000 cout=0 sum=01100011
* bcd_in1=00110101 bcd_in2=00101001 cout=0 sum=01100100
* bcd_in1=00110101 bcd_in2=00110000 cout=0 sum=01100101
* bcd_in1=00110101 bcd_in2=00110001 cout=0 sum=01100110
* bcd_in1=00110101 bcd_in2=00110010 cout=0 sum=01100111
* bcd_in1=00110101 bcd_in2=00110011 cout=0 sum=01101000
* bcd_in1=00110101 bcd_in2=00110100 cout=0 sum=01101001
* bcd_in1=00110101 bcd_in2=00110101 cout=0 sum=01110000
* bcd_in1=00110101 bcd_in2=00110110 cout=0 sum=01110001
* bcd_in1=00110101 bcd_in2=00110111 cout=0 sum=01110010
* bcd_in1=00110101 bcd_in2=00111000 cout=0 sum=01110011
* bcd_in1=00110101 bcd_in2=00111001 cout=0 sum=01110100
* bcd_in1=00110101 bcd_in2=01000000 cout=0 sum=01110101
* bcd_in1=00110101 bcd_in2=01000001 cout=0 sum=01110110
* bcd_in1=00110101 bcd_in2=01000010 cout=0 sum=01110111
* bcd_in1=00110101 bcd_in2=01000011 cout=0 sum=01111000
* bcd_in1=00110101 bcd_in2=01000100 cout=0 sum=01111001
* bcd_in1=00110101 bcd_in2=01000101 cout=0 sum=10000000
* bcd_in1=00110101 bcd_in2=01000110 cout=0 sum=10000001
* bcd_in1=00110101 bcd_in2=01000111 cout=0 sum=10000010
* bcd_in1=00110101 bcd_in2=01001000 cout=0 sum=10000011
* bcd_in1=00110101 bcd_in2=01001001 cout=0 sum=10000100
* bcd_in1=00110101 bcd_in2=01010000 cout=0 sum=10000101
* bcd_in1=00110101 bcd_in2=01010001 cout=0 sum=10000110
* bcd_in1=00110101 bcd_in2=01010010 cout=0 sum=10000111
* bcd_in1=00110101 bcd_in2=01010011 cout=0 sum=10001000
* bcd_in1=00110101 bcd_in2=01010100 cout=0 sum=10001001
* bcd_in1=00110101 bcd_in2=01010101 cout=0 sum=10010000
* bcd_in1=00110101 bcd_in2=01010110 cout=0 sum=10010001
* bcd_in1=00110101 bcd_in2=01010111 cout=0 sum=10010010
* bcd_in1=00110101 bcd_in2=01011000 cout=0 sum=10010011
* bcd_in1=00110101 bcd_in2=01011001 cout=0 sum=10010100
* bcd_in1=00110101 bcd_in2=01100000 cout=0 sum=10010101
* bcd_in1=00110101 bcd_in2=01100001 cout=0 sum=10010110
* bcd_in1=00110101 bcd_in2=01100010 cout=0 sum=10010111
* bcd_in1=00110101 bcd_in2=01100011 cout=0 sum=10011000
* bcd_in1=00110101 bcd_in2=01100100 cout=0 sum=10011001
* bcd_in1=00110101 bcd_in2=01100101 cout=1 sum=00000000
* bcd_in1=00110101 bcd_in2=01100110 cout=1 sum=00000001
* bcd_in1=00110101 bcd_in2=01100111 cout=1 sum=00000010
* bcd_in1=00110101 bcd_in2=01101000 cout=1 sum=00000011
* bcd_in1=00110101 bcd_in2=01101001 cout=1 sum=00000100
* bcd_in1=00110101 bcd_in2=01110000 cout=1 sum=00000101
* bcd_in1=00110101 bcd_in2=01110001 cout=1 sum=00000110
* bcd_in1=00110101 bcd_in2=01110010 cout=1 sum=00000111
* bcd_in1=00110101 bcd_in2=01110011 cout=1 sum=00001000
* bcd_in1=00110101 bcd_in2=01110100 cout=1 sum=00001001
* bcd_in1=00110101 bcd_in2=01110101 cout=1 sum=00010000
* bcd_in1=00110101 bcd_in2=01110110 cout=1 sum=00010001
* bcd_in1=00110101 bcd_in2=01110111 cout=1 sum=00010010
* bcd_in1=00110101 bcd_in2=01111000 cout=1 sum=00010011
* bcd_in1=00110101 bcd_in2=01111001 cout=1 sum=00010100
* bcd_in1=00110101 bcd_in2=10000000 cout=1 sum=00010101
* bcd_in1=00110101 bcd_in2=10000001 cout=1 sum=00010110
* bcd_in1=00110101 bcd_in2=10000010 cout=1 sum=00010111
* bcd_in1=00110101 bcd_in2=10000011 cout=1 sum=00011000
* bcd_in1=00110101 bcd_in2=10000100 cout=1 sum=00011001
* bcd_in1=00110101 bcd_in2=10000101 cout=1 sum=00100000
* bcd_in1=00110101 bcd_in2=10000110 cout=1 sum=00100001
* bcd_in1=00110101 bcd_in2=10000111 cout=1 sum=00100010
* bcd_in1=00110101 bcd_in2=10001000 cout=1 sum=00100011
* bcd_in1=00110101 bcd_in2=10001001 cout=1 sum=00100100
* bcd_in1=00110101 bcd_in2=10010000 cout=1 sum=00100101
* bcd_in1=00110101 bcd_in2=10010001 cout=1 sum=00100110
* bcd_in1=00110101 bcd_in2=10010010 cout=1 sum=00100111
* bcd_in1=00110101 bcd_in2=10010011 cout=1 sum=00101000
* bcd_in1=00110101 bcd_in2=10010100 cout=1 sum=00101001
* bcd_in1=00110101 bcd_in2=10010101 cout=1 sum=00110000
* bcd_in1=00110101 bcd_in2=10010110 cout=1 sum=00110001
* bcd_in1=00110101 bcd_in2=10010111 cout=1 sum=00110010
* bcd_in1=00110101 bcd_in2=10011000 cout=1 sum=00110011
* bcd_in1=00110101 bcd_in2=10011001 cout=1 sum=00110100
* bcd_in1=00110110 bcd_in2=00000000 cout=0 sum=00110110
* bcd_in1=00110110 bcd_in2=00000001 cout=0 sum=00110111
* bcd_in1=00110110 bcd_in2=00000010 cout=0 sum=00111000
* bcd_in1=00110110 bcd_in2=00000011 cout=0 sum=00111001
* bcd_in1=00110110 bcd_in2=00000100 cout=0 sum=01000000
* bcd_in1=00110110 bcd_in2=00000101 cout=0 sum=01000001
* bcd_in1=00110110 bcd_in2=00000110 cout=0 sum=01000010
* bcd_in1=00110110 bcd_in2=00000111 cout=0 sum=01000011
* bcd_in1=00110110 bcd_in2=00001000 cout=0 sum=01000100
* bcd_in1=00110110 bcd_in2=00001001 cout=0 sum=01000101
* bcd_in1=00110110 bcd_in2=00010000 cout=0 sum=01000110
* bcd_in1=00110110 bcd_in2=00010001 cout=0 sum=01000111
* bcd_in1=00110110 bcd_in2=00010010 cout=0 sum=01001000
* bcd_in1=00110110 bcd_in2=00010011 cout=0 sum=01001001
* bcd_in1=00110110 bcd_in2=00010100 cout=0 sum=01010000
* bcd_in1=00110110 bcd_in2=00010101 cout=0 sum=01010001
* bcd_in1=00110110 bcd_in2=00010110 cout=0 sum=01010010
* bcd_in1=00110110 bcd_in2=00010111 cout=0 sum=01010011
* bcd_in1=00110110 bcd_in2=00011000 cout=0 sum=01010100
* bcd_in1=00110110 bcd_in2=00011001 cout=0 sum=01010101
* bcd_in1=00110110 bcd_in2=00100000 cout=0 sum=01010110
* bcd_in1=00110110 bcd_in2=00100001 cout=0 sum=01010111
* bcd_in1=00110110 bcd_in2=00100010 cout=0 sum=01011000
* bcd_in1=00110110 bcd_in2=00100011 cout=0 sum=01011001
* bcd_in1=00110110 bcd_in2=00100100 cout=0 sum=01100000
* bcd_in1=00110110 bcd_in2=00100101 cout=0 sum=01100001
* bcd_in1=00110110 bcd_in2=00100110 cout=0 sum=01100010
* bcd_in1=00110110 bcd_in2=00100111 cout=0 sum=01100011
* bcd_in1=00110110 bcd_in2=00101000 cout=0 sum=01100100
* bcd_in1=00110110 bcd_in2=00101001 cout=0 sum=01100101
* bcd_in1=00110110 bcd_in2=00110000 cout=0 sum=01100110
* bcd_in1=00110110 bcd_in2=00110001 cout=0 sum=01100111
* bcd_in1=00110110 bcd_in2=00110010 cout=0 sum=01101000
* bcd_in1=00110110 bcd_in2=00110011 cout=0 sum=01101001
* bcd_in1=00110110 bcd_in2=00110100 cout=0 sum=01110000
* bcd_in1=00110110 bcd_in2=00110101 cout=0 sum=01110001
* bcd_in1=00110110 bcd_in2=00110110 cout=0 sum=01110010
* bcd_in1=00110110 bcd_in2=00110111 cout=0 sum=01110011
* bcd_in1=00110110 bcd_in2=00111000 cout=0 sum=01110100
* bcd_in1=00110110 bcd_in2=00111001 cout=0 sum=01110101
* bcd_in1=00110110 bcd_in2=01000000 cout=0 sum=01110110
* bcd_in1=00110110 bcd_in2=01000001 cout=0 sum=01110111
* bcd_in1=00110110 bcd_in2=01000010 cout=0 sum=01111000
* bcd_in1=00110110 bcd_in2=01000011 cout=0 sum=01111001
* bcd_in1=00110110 bcd_in2=01000100 cout=0 sum=10000000
* bcd_in1=00110110 bcd_in2=01000101 cout=0 sum=10000001
* bcd_in1=00110110 bcd_in2=01000110 cout=0 sum=10000010
* bcd_in1=00110110 bcd_in2=01000111 cout=0 sum=10000011
* bcd_in1=00110110 bcd_in2=01001000 cout=0 sum=10000100
* bcd_in1=00110110 bcd_in2=01001001 cout=0 sum=10000101
* bcd_in1=00110110 bcd_in2=01010000 cout=0 sum=10000110
* bcd_in1=00110110 bcd_in2=01010001 cout=0 sum=10000111
* bcd_in1=00110110 bcd_in2=01010010 cout=0 sum=10001000
* bcd_in1=00110110 bcd_in2=01010011 cout=0 sum=10001001
* bcd_in1=00110110 bcd_in2=01010100 cout=0 sum=10010000
* bcd_in1=00110110 bcd_in2=01010101 cout=0 sum=10010001
* bcd_in1=00110110 bcd_in2=01010110 cout=0 sum=10010010
* bcd_in1=00110110 bcd_in2=01010111 cout=0 sum=10010011
* bcd_in1=00110110 bcd_in2=01011000 cout=0 sum=10010100
* bcd_in1=00110110 bcd_in2=01011001 cout=0 sum=10010101
* bcd_in1=00110110 bcd_in2=01100000 cout=0 sum=10010110
* bcd_in1=00110110 bcd_in2=01100001 cout=0 sum=10010111
* bcd_in1=00110110 bcd_in2=01100010 cout=0 sum=10011000
* bcd_in1=00110110 bcd_in2=01100011 cout=0 sum=10011001
* bcd_in1=00110110 bcd_in2=01100100 cout=1 sum=00000000
* bcd_in1=00110110 bcd_in2=01100101 cout=1 sum=00000001
* bcd_in1=00110110 bcd_in2=01100110 cout=1 sum=00000010
* bcd_in1=00110110 bcd_in2=01100111 cout=1 sum=00000011
* bcd_in1=00110110 bcd_in2=01101000 cout=1 sum=00000100
* bcd_in1=00110110 bcd_in2=01101001 cout=1 sum=00000101
* bcd_in1=00110110 bcd_in2=01110000 cout=1 sum=00000110
* bcd_in1=00110110 bcd_in2=01110001 cout=1 sum=00000111
* bcd_in1=00110110 bcd_in2=01110010 cout=1 sum=00001000
* bcd_in1=00110110 bcd_in2=01110011 cout=1 sum=00001001
* bcd_in1=00110110 bcd_in2=01110100 cout=1 sum=00010000
* bcd_in1=00110110 bcd_in2=01110101 cout=1 sum=00010001
* bcd_in1=00110110 bcd_in2=01110110 cout=1 sum=00010010
* bcd_in1=00110110 bcd_in2=01110111 cout=1 sum=00010011
* bcd_in1=00110110 bcd_in2=01111000 cout=1 sum=00010100
* bcd_in1=00110110 bcd_in2=01111001 cout=1 sum=00010101
* bcd_in1=00110110 bcd_in2=10000000 cout=1 sum=00010110
* bcd_in1=00110110 bcd_in2=10000001 cout=1 sum=00010111
* bcd_in1=00110110 bcd_in2=10000010 cout=1 sum=00011000
* bcd_in1=00110110 bcd_in2=10000011 cout=1 sum=00011001
* bcd_in1=00110110 bcd_in2=10000100 cout=1 sum=00100000
* bcd_in1=00110110 bcd_in2=10000101 cout=1 sum=00100001
* bcd_in1=00110110 bcd_in2=10000110 cout=1 sum=00100010
* bcd_in1=00110110 bcd_in2=10000111 cout=1 sum=00100011
* bcd_in1=00110110 bcd_in2=10001000 cout=1 sum=00100100
* bcd_in1=00110110 bcd_in2=10001001 cout=1 sum=00100101
* bcd_in1=00110110 bcd_in2=10010000 cout=1 sum=00100110
* bcd_in1=00110110 bcd_in2=10010001 cout=1 sum=00100111
* bcd_in1=00110110 bcd_in2=10010010 cout=1 sum=00101000
* bcd_in1=00110110 bcd_in2=10010011 cout=1 sum=00101001
* bcd_in1=00110110 bcd_in2=10010100 cout=1 sum=00110000
* bcd_in1=00110110 bcd_in2=10010101 cout=1 sum=00110001
* bcd_in1=00110110 bcd_in2=10010110 cout=1 sum=00110010
* bcd_in1=00110110 bcd_in2=10010111 cout=1 sum=00110011
* bcd_in1=00110110 bcd_in2=10011000 cout=1 sum=00110100
* bcd_in1=00110110 bcd_in2=10011001 cout=1 sum=00110101
* bcd_in1=00110111 bcd_in2=00000000 cout=0 sum=00110111
* bcd_in1=00110111 bcd_in2=00000001 cout=0 sum=00111000
* bcd_in1=00110111 bcd_in2=00000010 cout=0 sum=00111001
* bcd_in1=00110111 bcd_in2=00000011 cout=0 sum=01000000
* bcd_in1=00110111 bcd_in2=00000100 cout=0 sum=01000001
* bcd_in1=00110111 bcd_in2=00000101 cout=0 sum=01000010
* bcd_in1=00110111 bcd_in2=00000110 cout=0 sum=01000011
* bcd_in1=00110111 bcd_in2=00000111 cout=0 sum=01000100
* bcd_in1=00110111 bcd_in2=00001000 cout=0 sum=01000101
* bcd_in1=00110111 bcd_in2=00001001 cout=0 sum=01000110
* bcd_in1=00110111 bcd_in2=00010000 cout=0 sum=01000111
* bcd_in1=00110111 bcd_in2=00010001 cout=0 sum=01001000
* bcd_in1=00110111 bcd_in2=00010010 cout=0 sum=01001001
* bcd_in1=00110111 bcd_in2=00010011 cout=0 sum=01010000
* bcd_in1=00110111 bcd_in2=00010100 cout=0 sum=01010001
* bcd_in1=00110111 bcd_in2=00010101 cout=0 sum=01010010
* bcd_in1=00110111 bcd_in2=00010110 cout=0 sum=01010011
* bcd_in1=00110111 bcd_in2=00010111 cout=0 sum=01010100
* bcd_in1=00110111 bcd_in2=00011000 cout=0 sum=01010101
* bcd_in1=00110111 bcd_in2=00011001 cout=0 sum=01010110
* bcd_in1=00110111 bcd_in2=00100000 cout=0 sum=01010111
* bcd_in1=00110111 bcd_in2=00100001 cout=0 sum=01011000
* bcd_in1=00110111 bcd_in2=00100010 cout=0 sum=01011001
* bcd_in1=00110111 bcd_in2=00100011 cout=0 sum=01100000
* bcd_in1=00110111 bcd_in2=00100100 cout=0 sum=01100001
* bcd_in1=00110111 bcd_in2=00100101 cout=0 sum=01100010
* bcd_in1=00110111 bcd_in2=00100110 cout=0 sum=01100011
* bcd_in1=00110111 bcd_in2=00100111 cout=0 sum=01100100
* bcd_in1=00110111 bcd_in2=00101000 cout=0 sum=01100101
* bcd_in1=00110111 bcd_in2=00101001 cout=0 sum=01100110
* bcd_in1=00110111 bcd_in2=00110000 cout=0 sum=01100111
* bcd_in1=00110111 bcd_in2=00110001 cout=0 sum=01101000
* bcd_in1=00110111 bcd_in2=00110010 cout=0 sum=01101001
* bcd_in1=00110111 bcd_in2=00110011 cout=0 sum=01110000
* bcd_in1=00110111 bcd_in2=00110100 cout=0 sum=01110001
* bcd_in1=00110111 bcd_in2=00110101 cout=0 sum=01110010
* bcd_in1=00110111 bcd_in2=00110110 cout=0 sum=01110011
* bcd_in1=00110111 bcd_in2=00110111 cout=0 sum=01110100
* bcd_in1=00110111 bcd_in2=00111000 cout=0 sum=01110101
* bcd_in1=00110111 bcd_in2=00111001 cout=0 sum=01110110
* bcd_in1=00110111 bcd_in2=01000000 cout=0 sum=01110111
* bcd_in1=00110111 bcd_in2=01000001 cout=0 sum=01111000
* bcd_in1=00110111 bcd_in2=01000010 cout=0 sum=01111001
* bcd_in1=00110111 bcd_in2=01000011 cout=0 sum=10000000
* bcd_in1=00110111 bcd_in2=01000100 cout=0 sum=10000001
* bcd_in1=00110111 bcd_in2=01000101 cout=0 sum=10000010
* bcd_in1=00110111 bcd_in2=01000110 cout=0 sum=10000011
* bcd_in1=00110111 bcd_in2=01000111 cout=0 sum=10000100
* bcd_in1=00110111 bcd_in2=01001000 cout=0 sum=10000101
* bcd_in1=00110111 bcd_in2=01001001 cout=0 sum=10000110
* bcd_in1=00110111 bcd_in2=01010000 cout=0 sum=10000111
* bcd_in1=00110111 bcd_in2=01010001 cout=0 sum=10001000
* bcd_in1=00110111 bcd_in2=01010010 cout=0 sum=10001001
* bcd_in1=00110111 bcd_in2=01010011 cout=0 sum=10010000
* bcd_in1=00110111 bcd_in2=01010100 cout=0 sum=10010001
* bcd_in1=00110111 bcd_in2=01010101 cout=0 sum=10010010
* bcd_in1=00110111 bcd_in2=01010110 cout=0 sum=10010011
* bcd_in1=00110111 bcd_in2=01010111 cout=0 sum=10010100
* bcd_in1=00110111 bcd_in2=01011000 cout=0 sum=10010101
* bcd_in1=00110111 bcd_in2=01011001 cout=0 sum=10010110
* bcd_in1=00110111 bcd_in2=01100000 cout=0 sum=10010111
* bcd_in1=00110111 bcd_in2=01100001 cout=0 sum=10011000
* bcd_in1=00110111 bcd_in2=01100010 cout=0 sum=10011001
* bcd_in1=00110111 bcd_in2=01100011 cout=1 sum=00000000
* bcd_in1=00110111 bcd_in2=01100100 cout=1 sum=00000001
* bcd_in1=00110111 bcd_in2=01100101 cout=1 sum=00000010
* bcd_in1=00110111 bcd_in2=01100110 cout=1 sum=00000011
* bcd_in1=00110111 bcd_in2=01100111 cout=1 sum=00000100
* bcd_in1=00110111 bcd_in2=01101000 cout=1 sum=00000101
* bcd_in1=00110111 bcd_in2=01101001 cout=1 sum=00000110
* bcd_in1=00110111 bcd_in2=01110000 cout=1 sum=00000111
* bcd_in1=00110111 bcd_in2=01110001 cout=1 sum=00001000
* bcd_in1=00110111 bcd_in2=01110010 cout=1 sum=00001001
* bcd_in1=00110111 bcd_in2=01110011 cout=1 sum=00010000
* bcd_in1=00110111 bcd_in2=01110100 cout=1 sum=00010001
* bcd_in1=00110111 bcd_in2=01110101 cout=1 sum=00010010
* bcd_in1=00110111 bcd_in2=01110110 cout=1 sum=00010011
* bcd_in1=00110111 bcd_in2=01110111 cout=1 sum=00010100
* bcd_in1=00110111 bcd_in2=01111000 cout=1 sum=00010101
* bcd_in1=00110111 bcd_in2=01111001 cout=1 sum=00010110
* bcd_in1=00110111 bcd_in2=10000000 cout=1 sum=00010111
* bcd_in1=00110111 bcd_in2=10000001 cout=1 sum=00011000
* bcd_in1=00110111 bcd_in2=10000010 cout=1 sum=00011001
* bcd_in1=00110111 bcd_in2=10000011 cout=1 sum=00100000
* bcd_in1=00110111 bcd_in2=10000100 cout=1 sum=00100001
* bcd_in1=00110111 bcd_in2=10000101 cout=1 sum=00100010
* bcd_in1=00110111 bcd_in2=10000110 cout=1 sum=00100011
* bcd_in1=00110111 bcd_in2=10000111 cout=1 sum=00100100
* bcd_in1=00110111 bcd_in2=10001000 cout=1 sum=00100101
* bcd_in1=00110111 bcd_in2=10001001 cout=1 sum=00100110
* bcd_in1=00110111 bcd_in2=10010000 cout=1 sum=00100111
* bcd_in1=00110111 bcd_in2=10010001 cout=1 sum=00101000
* bcd_in1=00110111 bcd_in2=10010010 cout=1 sum=00101001
* bcd_in1=00110111 bcd_in2=10010011 cout=1 sum=00110000
* bcd_in1=00110111 bcd_in2=10010100 cout=1 sum=00110001
* bcd_in1=00110111 bcd_in2=10010101 cout=1 sum=00110010
* bcd_in1=00110111 bcd_in2=10010110 cout=1 sum=00110011
* bcd_in1=00110111 bcd_in2=10010111 cout=1 sum=00110100
* bcd_in1=00110111 bcd_in2=10011000 cout=1 sum=00110101
* bcd_in1=00110111 bcd_in2=10011001 cout=1 sum=00110110
* bcd_in1=00111000 bcd_in2=00000000 cout=0 sum=00111000
* bcd_in1=00111000 bcd_in2=00000001 cout=0 sum=00111001
* bcd_in1=00111000 bcd_in2=00000010 cout=0 sum=01000000
* bcd_in1=00111000 bcd_in2=00000011 cout=0 sum=01000001
* bcd_in1=00111000 bcd_in2=00000100 cout=0 sum=01000010
* bcd_in1=00111000 bcd_in2=00000101 cout=0 sum=01000011
* bcd_in1=00111000 bcd_in2=00000110 cout=0 sum=01000100
* bcd_in1=00111000 bcd_in2=00000111 cout=0 sum=01000101
* bcd_in1=00111000 bcd_in2=00001000 cout=0 sum=01000110
* bcd_in1=00111000 bcd_in2=00001001 cout=0 sum=01000111
* bcd_in1=00111000 bcd_in2=00010000 cout=0 sum=01001000
* bcd_in1=00111000 bcd_in2=00010001 cout=0 sum=01001001
* bcd_in1=00111000 bcd_in2=00010010 cout=0 sum=01010000
* bcd_in1=00111000 bcd_in2=00010011 cout=0 sum=01010001
* bcd_in1=00111000 bcd_in2=00010100 cout=0 sum=01010010
* bcd_in1=00111000 bcd_in2=00010101 cout=0 sum=01010011
* bcd_in1=00111000 bcd_in2=00010110 cout=0 sum=01010100
* bcd_in1=00111000 bcd_in2=00010111 cout=0 sum=01010101
* bcd_in1=00111000 bcd_in2=00011000 cout=0 sum=01010110
* bcd_in1=00111000 bcd_in2=00011001 cout=0 sum=01010111
* bcd_in1=00111000 bcd_in2=00100000 cout=0 sum=01011000
* bcd_in1=00111000 bcd_in2=00100001 cout=0 sum=01011001
* bcd_in1=00111000 bcd_in2=00100010 cout=0 sum=01100000
* bcd_in1=00111000 bcd_in2=00100011 cout=0 sum=01100001
* bcd_in1=00111000 bcd_in2=00100100 cout=0 sum=01100010
* bcd_in1=00111000 bcd_in2=00100101 cout=0 sum=01100011
* bcd_in1=00111000 bcd_in2=00100110 cout=0 sum=01100100
* bcd_in1=00111000 bcd_in2=00100111 cout=0 sum=01100101
* bcd_in1=00111000 bcd_in2=00101000 cout=0 sum=01100110
* bcd_in1=00111000 bcd_in2=00101001 cout=0 sum=01100111
* bcd_in1=00111000 bcd_in2=00110000 cout=0 sum=01101000
* bcd_in1=00111000 bcd_in2=00110001 cout=0 sum=01101001
* bcd_in1=00111000 bcd_in2=00110010 cout=0 sum=01110000
* bcd_in1=00111000 bcd_in2=00110011 cout=0 sum=01110001
* bcd_in1=00111000 bcd_in2=00110100 cout=0 sum=01110010
* bcd_in1=00111000 bcd_in2=00110101 cout=0 sum=01110011
* bcd_in1=00111000 bcd_in2=00110110 cout=0 sum=01110100
* bcd_in1=00111000 bcd_in2=00110111 cout=0 sum=01110101
* bcd_in1=00111000 bcd_in2=00111000 cout=0 sum=01110110
* bcd_in1=00111000 bcd_in2=00111001 cout=0 sum=01110111
* bcd_in1=00111000 bcd_in2=01000000 cout=0 sum=01111000
* bcd_in1=00111000 bcd_in2=01000001 cout=0 sum=01111001
* bcd_in1=00111000 bcd_in2=01000010 cout=0 sum=10000000
* bcd_in1=00111000 bcd_in2=01000011 cout=0 sum=10000001
* bcd_in1=00111000 bcd_in2=01000100 cout=0 sum=10000010
* bcd_in1=00111000 bcd_in2=01000101 cout=0 sum=10000011
* bcd_in1=00111000 bcd_in2=01000110 cout=0 sum=10000100
* bcd_in1=00111000 bcd_in2=01000111 cout=0 sum=10000101
* bcd_in1=00111000 bcd_in2=01001000 cout=0 sum=10000110
* bcd_in1=00111000 bcd_in2=01001001 cout=0 sum=10000111
* bcd_in1=00111000 bcd_in2=01010000 cout=0 sum=10001000
* bcd_in1=00111000 bcd_in2=01010001 cout=0 sum=10001001
* bcd_in1=00111000 bcd_in2=01010010 cout=0 sum=10010000
* bcd_in1=00111000 bcd_in2=01010011 cout=0 sum=10010001
* bcd_in1=00111000 bcd_in2=01010100 cout=0 sum=10010010
* bcd_in1=00111000 bcd_in2=01010101 cout=0 sum=10010011
* bcd_in1=00111000 bcd_in2=01010110 cout=0 sum=10010100
* bcd_in1=00111000 bcd_in2=01010111 cout=0 sum=10010101
* bcd_in1=00111000 bcd_in2=01011000 cout=0 sum=10010110
* bcd_in1=00111000 bcd_in2=01011001 cout=0 sum=10010111
* bcd_in1=00111000 bcd_in2=01100000 cout=0 sum=10011000
* bcd_in1=00111000 bcd_in2=01100001 cout=0 sum=10011001
* bcd_in1=00111000 bcd_in2=01100010 cout=1 sum=00000000
* bcd_in1=00111000 bcd_in2=01100011 cout=1 sum=00000001
* bcd_in1=00111000 bcd_in2=01100100 cout=1 sum=00000010
* bcd_in1=00111000 bcd_in2=01100101 cout=1 sum=00000011
* bcd_in1=00111000 bcd_in2=01100110 cout=1 sum=00000100
* bcd_in1=00111000 bcd_in2=01100111 cout=1 sum=00000101
* bcd_in1=00111000 bcd_in2=01101000 cout=1 sum=00000110
* bcd_in1=00111000 bcd_in2=01101001 cout=1 sum=00000111
* bcd_in1=00111000 bcd_in2=01110000 cout=1 sum=00001000
* bcd_in1=00111000 bcd_in2=01110001 cout=1 sum=00001001
* bcd_in1=00111000 bcd_in2=01110010 cout=1 sum=00010000
* bcd_in1=00111000 bcd_in2=01110011 cout=1 sum=00010001
* bcd_in1=00111000 bcd_in2=01110100 cout=1 sum=00010010
* bcd_in1=00111000 bcd_in2=01110101 cout=1 sum=00010011
* bcd_in1=00111000 bcd_in2=01110110 cout=1 sum=00010100
* bcd_in1=00111000 bcd_in2=01110111 cout=1 sum=00010101
* bcd_in1=00111000 bcd_in2=01111000 cout=1 sum=00010110
* bcd_in1=00111000 bcd_in2=01111001 cout=1 sum=00010111
* bcd_in1=00111000 bcd_in2=10000000 cout=1 sum=00011000
* bcd_in1=00111000 bcd_in2=10000001 cout=1 sum=00011001
* bcd_in1=00111000 bcd_in2=10000010 cout=1 sum=00100000
* bcd_in1=00111000 bcd_in2=10000011 cout=1 sum=00100001
* bcd_in1=00111000 bcd_in2=10000100 cout=1 sum=00100010
* bcd_in1=00111000 bcd_in2=10000101 cout=1 sum=00100011
* bcd_in1=00111000 bcd_in2=10000110 cout=1 sum=00100100
* bcd_in1=00111000 bcd_in2=10000111 cout=1 sum=00100101
* bcd_in1=00111000 bcd_in2=10001000 cout=1 sum=00100110
* bcd_in1=00111000 bcd_in2=10001001 cout=1 sum=00100111
* bcd_in1=00111000 bcd_in2=10010000 cout=1 sum=00101000
* bcd_in1=00111000 bcd_in2=10010001 cout=1 sum=00101001
* bcd_in1=00111000 bcd_in2=10010010 cout=1 sum=00110000
* bcd_in1=00111000 bcd_in2=10010011 cout=1 sum=00110001
* bcd_in1=00111000 bcd_in2=10010100 cout=1 sum=00110010
* bcd_in1=00111000 bcd_in2=10010101 cout=1 sum=00110011
* bcd_in1=00111000 bcd_in2=10010110 cout=1 sum=00110100
* bcd_in1=00111000 bcd_in2=10010111 cout=1 sum=00110101
* bcd_in1=00111000 bcd_in2=10011000 cout=1 sum=00110110
* bcd_in1=00111000 bcd_in2=10011001 cout=1 sum=00110111
* bcd_in1=00111001 bcd_in2=00000000 cout=0 sum=00111001
* bcd_in1=00111001 bcd_in2=00000001 cout=0 sum=01000000
* bcd_in1=00111001 bcd_in2=00000010 cout=0 sum=01000001
* bcd_in1=00111001 bcd_in2=00000011 cout=0 sum=01000010
* bcd_in1=00111001 bcd_in2=00000100 cout=0 sum=01000011
* bcd_in1=00111001 bcd_in2=00000101 cout=0 sum=01000100
* bcd_in1=00111001 bcd_in2=00000110 cout=0 sum=01000101
* bcd_in1=00111001 bcd_in2=00000111 cout=0 sum=01000110
* bcd_in1=00111001 bcd_in2=00001000 cout=0 sum=01000111
* bcd_in1=00111001 bcd_in2=00001001 cout=0 sum=01001000
* bcd_in1=00111001 bcd_in2=00010000 cout=0 sum=01001001
* bcd_in1=00111001 bcd_in2=00010001 cout=0 sum=01010000
* bcd_in1=00111001 bcd_in2=00010010 cout=0 sum=01010001
* bcd_in1=00111001 bcd_in2=00010011 cout=0 sum=01010010
* bcd_in1=00111001 bcd_in2=00010100 cout=0 sum=01010011
* bcd_in1=00111001 bcd_in2=00010101 cout=0 sum=01010100
* bcd_in1=00111001 bcd_in2=00010110 cout=0 sum=01010101
* bcd_in1=00111001 bcd_in2=00010111 cout=0 sum=01010110
* bcd_in1=00111001 bcd_in2=00011000 cout=0 sum=01010111
* bcd_in1=00111001 bcd_in2=00011001 cout=0 sum=01011000
* bcd_in1=00111001 bcd_in2=00100000 cout=0 sum=01011001
* bcd_in1=00111001 bcd_in2=00100001 cout=0 sum=01100000
* bcd_in1=00111001 bcd_in2=00100010 cout=0 sum=01100001
* bcd_in1=00111001 bcd_in2=00100011 cout=0 sum=01100010
* bcd_in1=00111001 bcd_in2=00100100 cout=0 sum=01100011
* bcd_in1=00111001 bcd_in2=00100101 cout=0 sum=01100100
* bcd_in1=00111001 bcd_in2=00100110 cout=0 sum=01100101
* bcd_in1=00111001 bcd_in2=00100111 cout=0 sum=01100110
* bcd_in1=00111001 bcd_in2=00101000 cout=0 sum=01100111
* bcd_in1=00111001 bcd_in2=00101001 cout=0 sum=01101000
* bcd_in1=00111001 bcd_in2=00110000 cout=0 sum=01101001
* bcd_in1=00111001 bcd_in2=00110001 cout=0 sum=01110000
* bcd_in1=00111001 bcd_in2=00110010 cout=0 sum=01110001
* bcd_in1=00111001 bcd_in2=00110011 cout=0 sum=01110010
* bcd_in1=00111001 bcd_in2=00110100 cout=0 sum=01110011
* bcd_in1=00111001 bcd_in2=00110101 cout=0 sum=01110100
* bcd_in1=00111001 bcd_in2=00110110 cout=0 sum=01110101
* bcd_in1=00111001 bcd_in2=00110111 cout=0 sum=01110110
* bcd_in1=00111001 bcd_in2=00111000 cout=0 sum=01110111
* bcd_in1=00111001 bcd_in2=00111001 cout=0 sum=01111000
* bcd_in1=00111001 bcd_in2=01000000 cout=0 sum=01111001
* bcd_in1=00111001 bcd_in2=01000001 cout=0 sum=10000000
* bcd_in1=00111001 bcd_in2=01000010 cout=0 sum=10000001
* bcd_in1=00111001 bcd_in2=01000011 cout=0 sum=10000010
* bcd_in1=00111001 bcd_in2=01000100 cout=0 sum=10000011
* bcd_in1=00111001 bcd_in2=01000101 cout=0 sum=10000100
* bcd_in1=00111001 bcd_in2=01000110 cout=0 sum=10000101
* bcd_in1=00111001 bcd_in2=01000111 cout=0 sum=10000110
* bcd_in1=00111001 bcd_in2=01001000 cout=0 sum=10000111
* bcd_in1=00111001 bcd_in2=01001001 cout=0 sum=10001000
* bcd_in1=00111001 bcd_in2=01010000 cout=0 sum=10001001
* bcd_in1=00111001 bcd_in2=01010001 cout=0 sum=10010000
* bcd_in1=00111001 bcd_in2=01010010 cout=0 sum=10010001
* bcd_in1=00111001 bcd_in2=01010011 cout=0 sum=10010010
* bcd_in1=00111001 bcd_in2=01010100 cout=0 sum=10010011
* bcd_in1=00111001 bcd_in2=01010101 cout=0 sum=10010100
* bcd_in1=00111001 bcd_in2=01010110 cout=0 sum=10010101
* bcd_in1=00111001 bcd_in2=01010111 cout=0 sum=10010110
* bcd_in1=00111001 bcd_in2=01011000 cout=0 sum=10010111
* bcd_in1=00111001 bcd_in2=01011001 cout=0 sum=10011000
* bcd_in1=00111001 bcd_in2=01100000 cout=0 sum=10011001
* bcd_in1=00111001 bcd_in2=01100001 cout=1 sum=00000000
* bcd_in1=00111001 bcd_in2=01100010 cout=1 sum=00000001
* bcd_in1=00111001 bcd_in2=01100011 cout=1 sum=00000010
* bcd_in1=00111001 bcd_in2=01100100 cout=1 sum=00000011
* bcd_in1=00111001 bcd_in2=01100101 cout=1 sum=00000100
* bcd_in1=00111001 bcd_in2=01100110 cout=1 sum=00000101
* bcd_in1=00111001 bcd_in2=01100111 cout=1 sum=00000110
* bcd_in1=00111001 bcd_in2=01101000 cout=1 sum=00000111
* bcd_in1=00111001 bcd_in2=01101001 cout=1 sum=00001000
* bcd_in1=00111001 bcd_in2=01110000 cout=1 sum=00001001
* bcd_in1=00111001 bcd_in2=01110001 cout=1 sum=00010000
* bcd_in1=00111001 bcd_in2=01110010 cout=1 sum=00010001
* bcd_in1=00111001 bcd_in2=01110011 cout=1 sum=00010010
* bcd_in1=00111001 bcd_in2=01110100 cout=1 sum=00010011
* bcd_in1=00111001 bcd_in2=01110101 cout=1 sum=00010100
* bcd_in1=00111001 bcd_in2=01110110 cout=1 sum=00010101
* bcd_in1=00111001 bcd_in2=01110111 cout=1 sum=00010110
* bcd_in1=00111001 bcd_in2=01111000 cout=1 sum=00010111
* bcd_in1=00111001 bcd_in2=01111001 cout=1 sum=00011000
* bcd_in1=00111001 bcd_in2=10000000 cout=1 sum=00011001
* bcd_in1=00111001 bcd_in2=10000001 cout=1 sum=00100000
* bcd_in1=00111001 bcd_in2=10000010 cout=1 sum=00100001
* bcd_in1=00111001 bcd_in2=10000011 cout=1 sum=00100010
* bcd_in1=00111001 bcd_in2=10000100 cout=1 sum=00100011
* bcd_in1=00111001 bcd_in2=10000101 cout=1 sum=00100100
* bcd_in1=00111001 bcd_in2=10000110 cout=1 sum=00100101
* bcd_in1=00111001 bcd_in2=10000111 cout=1 sum=00100110
* bcd_in1=00111001 bcd_in2=10001000 cout=1 sum=00100111
* bcd_in1=00111001 bcd_in2=10001001 cout=1 sum=00101000
* bcd_in1=00111001 bcd_in2=10010000 cout=1 sum=00101001
* bcd_in1=00111001 bcd_in2=10010001 cout=1 sum=00110000
* bcd_in1=00111001 bcd_in2=10010010 cout=1 sum=00110001
* bcd_in1=00111001 bcd_in2=10010011 cout=1 sum=00110010
* bcd_in1=00111001 bcd_in2=10010100 cout=1 sum=00110011
* bcd_in1=00111001 bcd_in2=10010101 cout=1 sum=00110100
* bcd_in1=00111001 bcd_in2=10010110 cout=1 sum=00110101
* bcd_in1=00111001 bcd_in2=10010111 cout=1 sum=00110110
* bcd_in1=00111001 bcd_in2=10011000 cout=1 sum=00110111
* bcd_in1=00111001 bcd_in2=10011001 cout=1 sum=00111000
* bcd_in1=01000000 bcd_in2=00000000 cout=0 sum=01000000
* bcd_in1=01000000 bcd_in2=00000001 cout=0 sum=01000001
* bcd_in1=01000000 bcd_in2=00000010 cout=0 sum=01000010
* bcd_in1=01000000 bcd_in2=00000011 cout=0 sum=01000011
* bcd_in1=01000000 bcd_in2=00000100 cout=0 sum=01000100
* bcd_in1=01000000 bcd_in2=00000101 cout=0 sum=01000101
* bcd_in1=01000000 bcd_in2=00000110 cout=0 sum=01000110
* bcd_in1=01000000 bcd_in2=00000111 cout=0 sum=01000111
* bcd_in1=01000000 bcd_in2=00001000 cout=0 sum=01001000
* bcd_in1=01000000 bcd_in2=00001001 cout=0 sum=01001001
* bcd_in1=01000000 bcd_in2=00010000 cout=0 sum=01010000
* bcd_in1=01000000 bcd_in2=00010001 cout=0 sum=01010001
* bcd_in1=01000000 bcd_in2=00010010 cout=0 sum=01010010
* bcd_in1=01000000 bcd_in2=00010011 cout=0 sum=01010011
* bcd_in1=01000000 bcd_in2=00010100 cout=0 sum=01010100
* bcd_in1=01000000 bcd_in2=00010101 cout=0 sum=01010101
* bcd_in1=01000000 bcd_in2=00010110 cout=0 sum=01010110
* bcd_in1=01000000 bcd_in2=00010111 cout=0 sum=01010111
* bcd_in1=01000000 bcd_in2=00011000 cout=0 sum=01011000
* bcd_in1=01000000 bcd_in2=00011001 cout=0 sum=01011001
* bcd_in1=01000000 bcd_in2=00100000 cout=0 sum=01100000
* bcd_in1=01000000 bcd_in2=00100001 cout=0 sum=01100001
* bcd_in1=01000000 bcd_in2=00100010 cout=0 sum=01100010
* bcd_in1=01000000 bcd_in2=00100011 cout=0 sum=01100011
* bcd_in1=01000000 bcd_in2=00100100 cout=0 sum=01100100
* bcd_in1=01000000 bcd_in2=00100101 cout=0 sum=01100101
* bcd_in1=01000000 bcd_in2=00100110 cout=0 sum=01100110
* bcd_in1=01000000 bcd_in2=00100111 cout=0 sum=01100111
* bcd_in1=01000000 bcd_in2=00101000 cout=0 sum=01101000
* bcd_in1=01000000 bcd_in2=00101001 cout=0 sum=01101001
* bcd_in1=01000000 bcd_in2=00110000 cout=0 sum=01110000
* bcd_in1=01000000 bcd_in2=00110001 cout=0 sum=01110001
* bcd_in1=01000000 bcd_in2=00110010 cout=0 sum=01110010
* bcd_in1=01000000 bcd_in2=00110011 cout=0 sum=01110011
* bcd_in1=01000000 bcd_in2=00110100 cout=0 sum=01110100
* bcd_in1=01000000 bcd_in2=00110101 cout=0 sum=01110101
* bcd_in1=01000000 bcd_in2=00110110 cout=0 sum=01110110
* bcd_in1=01000000 bcd_in2=00110111 cout=0 sum=01110111
* bcd_in1=01000000 bcd_in2=00111000 cout=0 sum=01111000
* bcd_in1=01000000 bcd_in2=00111001 cout=0 sum=01111001
* bcd_in1=01000000 bcd_in2=01000000 cout=0 sum=10000000
* bcd_in1=01000000 bcd_in2=01000001 cout=0 sum=10000001
* bcd_in1=01000000 bcd_in2=01000010 cout=0 sum=10000010
* bcd_in1=01000000 bcd_in2=01000011 cout=0 sum=10000011
* bcd_in1=01000000 bcd_in2=01000100 cout=0 sum=10000100
* bcd_in1=01000000 bcd_in2=01000101 cout=0 sum=10000101
* bcd_in1=01000000 bcd_in2=01000110 cout=0 sum=10000110
* bcd_in1=01000000 bcd_in2=01000111 cout=0 sum=10000111
* bcd_in1=01000000 bcd_in2=01001000 cout=0 sum=10001000
* bcd_in1=01000000 bcd_in2=01001001 cout=0 sum=10001001
* bcd_in1=01000000 bcd_in2=01010000 cout=0 sum=10010000
* bcd_in1=01000000 bcd_in2=01010001 cout=0 sum=10010001
* bcd_in1=01000000 bcd_in2=01010010 cout=0 sum=10010010
* bcd_in1=01000000 bcd_in2=01010011 cout=0 sum=10010011
* bcd_in1=01000000 bcd_in2=01010100 cout=0 sum=10010100
* bcd_in1=01000000 bcd_in2=01010101 cout=0 sum=10010101
* bcd_in1=01000000 bcd_in2=01010110 cout=0 sum=10010110
* bcd_in1=01000000 bcd_in2=01010111 cout=0 sum=10010111
* bcd_in1=01000000 bcd_in2=01011000 cout=0 sum=10011000
* bcd_in1=01000000 bcd_in2=01011001 cout=0 sum=10011001
* bcd_in1=01000000 bcd_in2=01100000 cout=1 sum=00000000
* bcd_in1=01000000 bcd_in2=01100001 cout=1 sum=00000001
* bcd_in1=01000000 bcd_in2=01100010 cout=1 sum=00000010
* bcd_in1=01000000 bcd_in2=01100011 cout=1 sum=00000011
* bcd_in1=01000000 bcd_in2=01100100 cout=1 sum=00000100
* bcd_in1=01000000 bcd_in2=01100101 cout=1 sum=00000101
* bcd_in1=01000000 bcd_in2=01100110 cout=1 sum=00000110
* bcd_in1=01000000 bcd_in2=01100111 cout=1 sum=00000111
* bcd_in1=01000000 bcd_in2=01101000 cout=1 sum=00001000
* bcd_in1=01000000 bcd_in2=01101001 cout=1 sum=00001001
* bcd_in1=01000000 bcd_in2=01110000 cout=1 sum=00010000
* bcd_in1=01000000 bcd_in2=01110001 cout=1 sum=00010001
* bcd_in1=01000000 bcd_in2=01110010 cout=1 sum=00010010
* bcd_in1=01000000 bcd_in2=01110011 cout=1 sum=00010011
* bcd_in1=01000000 bcd_in2=01110100 cout=1 sum=00010100
* bcd_in1=01000000 bcd_in2=01110101 cout=1 sum=00010101
* bcd_in1=01000000 bcd_in2=01110110 cout=1 sum=00010110
* bcd_in1=01000000 bcd_in2=01110111 cout=1 sum=00010111
* bcd_in1=01000000 bcd_in2=01111000 cout=1 sum=00011000
* bcd_in1=01000000 bcd_in2=01111001 cout=1 sum=00011001
* bcd_in1=01000000 bcd_in2=10000000 cout=1 sum=00100000
* bcd_in1=01000000 bcd_in2=10000001 cout=1 sum=00100001
* bcd_in1=01000000 bcd_in2=10000010 cout=1 sum=00100010
* bcd_in1=01000000 bcd_in2=10000011 cout=1 sum=00100011
* bcd_in1=01000000 bcd_in2=10000100 cout=1 sum=00100100
* bcd_in1=01000000 bcd_in2=10000101 cout=1 sum=00100101
* bcd_in1=01000000 bcd_in2=10000110 cout=1 sum=00100110
* bcd_in1=01000000 bcd_in2=10000111 cout=1 sum=00100111
* bcd_in1=01000000 bcd_in2=10001000 cout=1 sum=00101000
* bcd_in1=01000000 bcd_in2=10001001 cout=1 sum=00101001
* bcd_in1=01000000 bcd_in2=10010000 cout=1 sum=00110000
* bcd_in1=01000000 bcd_in2=10010001 cout=1 sum=00110001
* bcd_in1=01000000 bcd_in2=10010010 cout=1 sum=00110010
* bcd_in1=01000000 bcd_in2=10010011 cout=1 sum=00110011
* bcd_in1=01000000 bcd_in2=10010100 cout=1 sum=00110100
* bcd_in1=01000000 bcd_in2=10010101 cout=1 sum=00110101
* bcd_in1=01000000 bcd_in2=10010110 cout=1 sum=00110110
* bcd_in1=01000000 bcd_in2=10010111 cout=1 sum=00110111
* bcd_in1=01000000 bcd_in2=10011000 cout=1 sum=00111000
* bcd_in1=01000000 bcd_in2=10011001 cout=1 sum=00111001
* bcd_in1=01000001 bcd_in2=00000000 cout=0 sum=01000001
* bcd_in1=01000001 bcd_in2=00000001 cout=0 sum=01000010
* bcd_in1=01000001 bcd_in2=00000010 cout=0 sum=01000011
* bcd_in1=01000001 bcd_in2=00000011 cout=0 sum=01000100
* bcd_in1=01000001 bcd_in2=00000100 cout=0 sum=01000101
* bcd_in1=01000001 bcd_in2=00000101 cout=0 sum=01000110
* bcd_in1=01000001 bcd_in2=00000110 cout=0 sum=01000111
* bcd_in1=01000001 bcd_in2=00000111 cout=0 sum=01001000
* bcd_in1=01000001 bcd_in2=00001000 cout=0 sum=01001001
* bcd_in1=01000001 bcd_in2=00001001 cout=0 sum=01010000
* bcd_in1=01000001 bcd_in2=00010000 cout=0 sum=01010001
* bcd_in1=01000001 bcd_in2=00010001 cout=0 sum=01010010
* bcd_in1=01000001 bcd_in2=00010010 cout=0 sum=01010011
* bcd_in1=01000001 bcd_in2=00010011 cout=0 sum=01010100
* bcd_in1=01000001 bcd_in2=00010100 cout=0 sum=01010101
* bcd_in1=01000001 bcd_in2=00010101 cout=0 sum=01010110
* bcd_in1=01000001 bcd_in2=00010110 cout=0 sum=01010111
* bcd_in1=01000001 bcd_in2=00010111 cout=0 sum=01011000
* bcd_in1=01000001 bcd_in2=00011000 cout=0 sum=01011001
* bcd_in1=01000001 bcd_in2=00011001 cout=0 sum=01100000
* bcd_in1=01000001 bcd_in2=00100000 cout=0 sum=01100001
* bcd_in1=01000001 bcd_in2=00100001 cout=0 sum=01100010
* bcd_in1=01000001 bcd_in2=00100010 cout=0 sum=01100011
* bcd_in1=01000001 bcd_in2=00100011 cout=0 sum=01100100
* bcd_in1=01000001 bcd_in2=00100100 cout=0 sum=01100101
* bcd_in1=01000001 bcd_in2=00100101 cout=0 sum=01100110
* bcd_in1=01000001 bcd_in2=00100110 cout=0 sum=01100111
* bcd_in1=01000001 bcd_in2=00100111 cout=0 sum=01101000
* bcd_in1=01000001 bcd_in2=00101000 cout=0 sum=01101001
* bcd_in1=01000001 bcd_in2=00101001 cout=0 sum=01110000
* bcd_in1=01000001 bcd_in2=00110000 cout=0 sum=01110001
* bcd_in1=01000001 bcd_in2=00110001 cout=0 sum=01110010
* bcd_in1=01000001 bcd_in2=00110010 cout=0 sum=01110011
* bcd_in1=01000001 bcd_in2=00110011 cout=0 sum=01110100
* bcd_in1=01000001 bcd_in2=00110100 cout=0 sum=01110101
* bcd_in1=01000001 bcd_in2=00110101 cout=0 sum=01110110
* bcd_in1=01000001 bcd_in2=00110110 cout=0 sum=01110111
* bcd_in1=01000001 bcd_in2=00110111 cout=0 sum=01111000
* bcd_in1=01000001 bcd_in2=00111000 cout=0 sum=01111001
* bcd_in1=01000001 bcd_in2=00111001 cout=0 sum=10000000
* bcd_in1=01000001 bcd_in2=01000000 cout=0 sum=10000001
* bcd_in1=01000001 bcd_in2=01000001 cout=0 sum=10000010
* bcd_in1=01000001 bcd_in2=01000010 cout=0 sum=10000011
* bcd_in1=01000001 bcd_in2=01000011 cout=0 sum=10000100
* bcd_in1=01000001 bcd_in2=01000100 cout=0 sum=10000101
* bcd_in1=01000001 bcd_in2=01000101 cout=0 sum=10000110
* bcd_in1=01000001 bcd_in2=01000110 cout=0 sum=10000111
* bcd_in1=01000001 bcd_in2=01000111 cout=0 sum=10001000
* bcd_in1=01000001 bcd_in2=01001000 cout=0 sum=10001001
* bcd_in1=01000001 bcd_in2=01001001 cout=0 sum=10010000
* bcd_in1=01000001 bcd_in2=01010000 cout=0 sum=10010001
* bcd_in1=01000001 bcd_in2=01010001 cout=0 sum=10010010
* bcd_in1=01000001 bcd_in2=01010010 cout=0 sum=10010011
* bcd_in1=01000001 bcd_in2=01010011 cout=0 sum=10010100
* bcd_in1=01000001 bcd_in2=01010100 cout=0 sum=10010101
* bcd_in1=01000001 bcd_in2=01010101 cout=0 sum=10010110
* bcd_in1=01000001 bcd_in2=01010110 cout=0 sum=10010111
* bcd_in1=01000001 bcd_in2=01010111 cout=0 sum=10011000
* bcd_in1=01000001 bcd_in2=01011000 cout=0 sum=10011001
* bcd_in1=01000001 bcd_in2=01011001 cout=1 sum=00000000
* bcd_in1=01000001 bcd_in2=01100000 cout=1 sum=00000001
* bcd_in1=01000001 bcd_in2=01100001 cout=1 sum=00000010
* bcd_in1=01000001 bcd_in2=01100010 cout=1 sum=00000011
* bcd_in1=01000001 bcd_in2=01100011 cout=1 sum=00000100
* bcd_in1=01000001 bcd_in2=01100100 cout=1 sum=00000101
* bcd_in1=01000001 bcd_in2=01100101 cout=1 sum=00000110
* bcd_in1=01000001 bcd_in2=01100110 cout=1 sum=00000111
* bcd_in1=01000001 bcd_in2=01100111 cout=1 sum=00001000
* bcd_in1=01000001 bcd_in2=01101000 cout=1 sum=00001001
* bcd_in1=01000001 bcd_in2=01101001 cout=1 sum=00010000
* bcd_in1=01000001 bcd_in2=01110000 cout=1 sum=00010001
* bcd_in1=01000001 bcd_in2=01110001 cout=1 sum=00010010
* bcd_in1=01000001 bcd_in2=01110010 cout=1 sum=00010011
* bcd_in1=01000001 bcd_in2=01110011 cout=1 sum=00010100
* bcd_in1=01000001 bcd_in2=01110100 cout=1 sum=00010101
* bcd_in1=01000001 bcd_in2=01110101 cout=1 sum=00010110
* bcd_in1=01000001 bcd_in2=01110110 cout=1 sum=00010111
* bcd_in1=01000001 bcd_in2=01110111 cout=1 sum=00011000
* bcd_in1=01000001 bcd_in2=01111000 cout=1 sum=00011001
* bcd_in1=01000001 bcd_in2=01111001 cout=1 sum=00100000
* bcd_in1=01000001 bcd_in2=10000000 cout=1 sum=00100001
* bcd_in1=01000001 bcd_in2=10000001 cout=1 sum=00100010
* bcd_in1=01000001 bcd_in2=10000010 cout=1 sum=00100011
* bcd_in1=01000001 bcd_in2=10000011 cout=1 sum=00100100
* bcd_in1=01000001 bcd_in2=10000100 cout=1 sum=00100101
* bcd_in1=01000001 bcd_in2=10000101 cout=1 sum=00100110
* bcd_in1=01000001 bcd_in2=10000110 cout=1 sum=00100111
* bcd_in1=01000001 bcd_in2=10000111 cout=1 sum=00101000
* bcd_in1=01000001 bcd_in2=10001000 cout=1 sum=00101001
* bcd_in1=01000001 bcd_in2=10001001 cout=1 sum=00110000
* bcd_in1=01000001 bcd_in2=10010000 cout=1 sum=00110001
* bcd_in1=01000001 bcd_in2=10010001 cout=1 sum=00110010
* bcd_in1=01000001 bcd_in2=10010010 cout=1 sum=00110011
* bcd_in1=01000001 bcd_in2=10010011 cout=1 sum=00110100
* bcd_in1=01000001 bcd_in2=10010100 cout=1 sum=00110101
* bcd_in1=01000001 bcd_in2=10010101 cout=1 sum=00110110
* bcd_in1=01000001 bcd_in2=10010110 cout=1 sum=00110111
* bcd_in1=01000001 bcd_in2=10010111 cout=1 sum=00111000
* bcd_in1=01000001 bcd_in2=10011000 cout=1 sum=00111001
* bcd_in1=01000001 bcd_in2=10011001 cout=1 sum=01000000
* bcd_in1=01000010 bcd_in2=00000000 cout=0 sum=01000010
* bcd_in1=01000010 bcd_in2=00000001 cout=0 sum=01000011
* bcd_in1=01000010 bcd_in2=00000010 cout=0 sum=01000100
* bcd_in1=01000010 bcd_in2=00000011 cout=0 sum=01000101
* bcd_in1=01000010 bcd_in2=00000100 cout=0 sum=01000110
* bcd_in1=01000010 bcd_in2=00000101 cout=0 sum=01000111
* bcd_in1=01000010 bcd_in2=00000110 cout=0 sum=01001000
* bcd_in1=01000010 bcd_in2=00000111 cout=0 sum=01001001
* bcd_in1=01000010 bcd_in2=00001000 cout=0 sum=01010000
* bcd_in1=01000010 bcd_in2=00001001 cout=0 sum=01010001
* bcd_in1=01000010 bcd_in2=00010000 cout=0 sum=01010010
* bcd_in1=01000010 bcd_in2=00010001 cout=0 sum=01010011
* bcd_in1=01000010 bcd_in2=00010010 cout=0 sum=01010100
* bcd_in1=01000010 bcd_in2=00010011 cout=0 sum=01010101
* bcd_in1=01000010 bcd_in2=00010100 cout=0 sum=01010110
* bcd_in1=01000010 bcd_in2=00010101 cout=0 sum=01010111
* bcd_in1=01000010 bcd_in2=00010110 cout=0 sum=01011000
* bcd_in1=01000010 bcd_in2=00010111 cout=0 sum=01011001
* bcd_in1=01000010 bcd_in2=00011000 cout=0 sum=01100000
* bcd_in1=01000010 bcd_in2=00011001 cout=0 sum=01100001
* bcd_in1=01000010 bcd_in2=00100000 cout=0 sum=01100010
* bcd_in1=01000010 bcd_in2=00100001 cout=0 sum=01100011
* bcd_in1=01000010 bcd_in2=00100010 cout=0 sum=01100100
* bcd_in1=01000010 bcd_in2=00100011 cout=0 sum=01100101
* bcd_in1=01000010 bcd_in2=00100100 cout=0 sum=01100110
* bcd_in1=01000010 bcd_in2=00100101 cout=0 sum=01100111
* bcd_in1=01000010 bcd_in2=00100110 cout=0 sum=01101000
* bcd_in1=01000010 bcd_in2=00100111 cout=0 sum=01101001
* bcd_in1=01000010 bcd_in2=00101000 cout=0 sum=01110000
* bcd_in1=01000010 bcd_in2=00101001 cout=0 sum=01110001
* bcd_in1=01000010 bcd_in2=00110000 cout=0 sum=01110010
* bcd_in1=01000010 bcd_in2=00110001 cout=0 sum=01110011
* bcd_in1=01000010 bcd_in2=00110010 cout=0 sum=01110100
* bcd_in1=01000010 bcd_in2=00110011 cout=0 sum=01110101
* bcd_in1=01000010 bcd_in2=00110100 cout=0 sum=01110110
* bcd_in1=01000010 bcd_in2=00110101 cout=0 sum=01110111
* bcd_in1=01000010 bcd_in2=00110110 cout=0 sum=01111000
* bcd_in1=01000010 bcd_in2=00110111 cout=0 sum=01111001
* bcd_in1=01000010 bcd_in2=00111000 cout=0 sum=10000000
* bcd_in1=01000010 bcd_in2=00111001 cout=0 sum=10000001
* bcd_in1=01000010 bcd_in2=01000000 cout=0 sum=10000010
* bcd_in1=01000010 bcd_in2=01000001 cout=0 sum=10000011
* bcd_in1=01000010 bcd_in2=01000010 cout=0 sum=10000100
* bcd_in1=01000010 bcd_in2=01000011 cout=0 sum=10000101
* bcd_in1=01000010 bcd_in2=01000100 cout=0 sum=10000110
* bcd_in1=01000010 bcd_in2=01000101 cout=0 sum=10000111
* bcd_in1=01000010 bcd_in2=01000110 cout=0 sum=10001000
* bcd_in1=01000010 bcd_in2=01000111 cout=0 sum=10001001
* bcd_in1=01000010 bcd_in2=01001000 cout=0 sum=10010000
* bcd_in1=01000010 bcd_in2=01001001 cout=0 sum=10010001
* bcd_in1=01000010 bcd_in2=01010000 cout=0 sum=10010010
* bcd_in1=01000010 bcd_in2=01010001 cout=0 sum=10010011
* bcd_in1=01000010 bcd_in2=01010010 cout=0 sum=10010100
* bcd_in1=01000010 bcd_in2=01010011 cout=0 sum=10010101
* bcd_in1=01000010 bcd_in2=01010100 cout=0 sum=10010110
* bcd_in1=01000010 bcd_in2=01010101 cout=0 sum=10010111
* bcd_in1=01000010 bcd_in2=01010110 cout=0 sum=10011000
* bcd_in1=01000010 bcd_in2=01010111 cout=0 sum=10011001
* bcd_in1=01000010 bcd_in2=01011000 cout=1 sum=00000000
* bcd_in1=01000010 bcd_in2=01011001 cout=1 sum=00000001
* bcd_in1=01000010 bcd_in2=01100000 cout=1 sum=00000010
* bcd_in1=01000010 bcd_in2=01100001 cout=1 sum=00000011
* bcd_in1=01000010 bcd_in2=01100010 cout=1 sum=00000100
* bcd_in1=01000010 bcd_in2=01100011 cout=1 sum=00000101
* bcd_in1=01000010 bcd_in2=01100100 cout=1 sum=00000110
* bcd_in1=01000010 bcd_in2=01100101 cout=1 sum=00000111
* bcd_in1=01000010 bcd_in2=01100110 cout=1 sum=00001000
* bcd_in1=01000010 bcd_in2=01100111 cout=1 sum=00001001
* bcd_in1=01000010 bcd_in2=01101000 cout=1 sum=00010000
* bcd_in1=01000010 bcd_in2=01101001 cout=1 sum=00010001
* bcd_in1=01000010 bcd_in2=01110000 cout=1 sum=00010010
* bcd_in1=01000010 bcd_in2=01110001 cout=1 sum=00010011
* bcd_in1=01000010 bcd_in2=01110010 cout=1 sum=00010100
* bcd_in1=01000010 bcd_in2=01110011 cout=1 sum=00010101
* bcd_in1=01000010 bcd_in2=01110100 cout=1 sum=00010110
* bcd_in1=01000010 bcd_in2=01110101 cout=1 sum=00010111
* bcd_in1=01000010 bcd_in2=01110110 cout=1 sum=00011000
* bcd_in1=01000010 bcd_in2=01110111 cout=1 sum=00011001
* bcd_in1=01000010 bcd_in2=01111000 cout=1 sum=00100000
* bcd_in1=01000010 bcd_in2=01111001 cout=1 sum=00100001
* bcd_in1=01000010 bcd_in2=10000000 cout=1 sum=00100010
* bcd_in1=01000010 bcd_in2=10000001 cout=1 sum=00100011
* bcd_in1=01000010 bcd_in2=10000010 cout=1 sum=00100100
* bcd_in1=01000010 bcd_in2=10000011 cout=1 sum=00100101
* bcd_in1=01000010 bcd_in2=10000100 cout=1 sum=00100110
* bcd_in1=01000010 bcd_in2=10000101 cout=1 sum=00100111
* bcd_in1=01000010 bcd_in2=10000110 cout=1 sum=00101000
* bcd_in1=01000010 bcd_in2=10000111 cout=1 sum=00101001
* bcd_in1=01000010 bcd_in2=10001000 cout=1 sum=00110000
* bcd_in1=01000010 bcd_in2=10001001 cout=1 sum=00110001
* bcd_in1=01000010 bcd_in2=10010000 cout=1 sum=00110010
* bcd_in1=01000010 bcd_in2=10010001 cout=1 sum=00110011
* bcd_in1=01000010 bcd_in2=10010010 cout=1 sum=00110100
* bcd_in1=01000010 bcd_in2=10010011 cout=1 sum=00110101
* bcd_in1=01000010 bcd_in2=10010100 cout=1 sum=00110110
* bcd_in1=01000010 bcd_in2=10010101 cout=1 sum=00110111
* bcd_in1=01000010 bcd_in2=10010110 cout=1 sum=00111000
* bcd_in1=01000010 bcd_in2=10010111 cout=1 sum=00111001
* bcd_in1=01000010 bcd_in2=10011000 cout=1 sum=01000000
* bcd_in1=01000010 bcd_in2=10011001 cout=1 sum=01000001
* bcd_in1=01000011 bcd_in2=00000000 cout=0 sum=01000011
* bcd_in1=01000011 bcd_in2=00000001 cout=0 sum=01000100
* bcd_in1=01000011 bcd_in2=00000010 cout=0 sum=01000101
* bcd_in1=01000011 bcd_in2=00000011 cout=0 sum=01000110
* bcd_in1=01000011 bcd_in2=00000100 cout=0 sum=01000111
* bcd_in1=01000011 bcd_in2=00000101 cout=0 sum=01001000
* bcd_in1=01000011 bcd_in2=00000110 cout=0 sum=01001001
* bcd_in1=01000011 bcd_in2=00000111 cout=0 sum=01010000
* bcd_in1=01000011 bcd_in2=00001000 cout=0 sum=01010001
* bcd_in1=01000011 bcd_in2=00001001 cout=0 sum=01010010
* bcd_in1=01000011 bcd_in2=00010000 cout=0 sum=01010011
* bcd_in1=01000011 bcd_in2=00010001 cout=0 sum=01010100
* bcd_in1=01000011 bcd_in2=00010010 cout=0 sum=01010101
* bcd_in1=01000011 bcd_in2=00010011 cout=0 sum=01010110
* bcd_in1=01000011 bcd_in2=00010100 cout=0 sum=01010111
* bcd_in1=01000011 bcd_in2=00010101 cout=0 sum=01011000
* bcd_in1=01000011 bcd_in2=00010110 cout=0 sum=01011001
* bcd_in1=01000011 bcd_in2=00010111 cout=0 sum=01100000
* bcd_in1=01000011 bcd_in2=00011000 cout=0 sum=01100001
* bcd_in1=01000011 bcd_in2=00011001 cout=0 sum=01100010
* bcd_in1=01000011 bcd_in2=00100000 cout=0 sum=01100011
* bcd_in1=01000011 bcd_in2=00100001 cout=0 sum=01100100
* bcd_in1=01000011 bcd_in2=00100010 cout=0 sum=01100101
* bcd_in1=01000011 bcd_in2=00100011 cout=0 sum=01100110
* bcd_in1=01000011 bcd_in2=00100100 cout=0 sum=01100111
* bcd_in1=01000011 bcd_in2=00100101 cout=0 sum=01101000
* bcd_in1=01000011 bcd_in2=00100110 cout=0 sum=01101001
* bcd_in1=01000011 bcd_in2=00100111 cout=0 sum=01110000
* bcd_in1=01000011 bcd_in2=00101000 cout=0 sum=01110001
* bcd_in1=01000011 bcd_in2=00101001 cout=0 sum=01110010
* bcd_in1=01000011 bcd_in2=00110000 cout=0 sum=01110011
* bcd_in1=01000011 bcd_in2=00110001 cout=0 sum=01110100
* bcd_in1=01000011 bcd_in2=00110010 cout=0 sum=01110101
* bcd_in1=01000011 bcd_in2=00110011 cout=0 sum=01110110
* bcd_in1=01000011 bcd_in2=00110100 cout=0 sum=01110111
* bcd_in1=01000011 bcd_in2=00110101 cout=0 sum=01111000
* bcd_in1=01000011 bcd_in2=00110110 cout=0 sum=01111001
* bcd_in1=01000011 bcd_in2=00110111 cout=0 sum=10000000
* bcd_in1=01000011 bcd_in2=00111000 cout=0 sum=10000001
* bcd_in1=01000011 bcd_in2=00111001 cout=0 sum=10000010
* bcd_in1=01000011 bcd_in2=01000000 cout=0 sum=10000011
* bcd_in1=01000011 bcd_in2=01000001 cout=0 sum=10000100
* bcd_in1=01000011 bcd_in2=01000010 cout=0 sum=10000101
* bcd_in1=01000011 bcd_in2=01000011 cout=0 sum=10000110
* bcd_in1=01000011 bcd_in2=01000100 cout=0 sum=10000111
* bcd_in1=01000011 bcd_in2=01000101 cout=0 sum=10001000
* bcd_in1=01000011 bcd_in2=01000110 cout=0 sum=10001001
* bcd_in1=01000011 bcd_in2=01000111 cout=0 sum=10010000
* bcd_in1=01000011 bcd_in2=01001000 cout=0 sum=10010001
* bcd_in1=01000011 bcd_in2=01001001 cout=0 sum=10010010
* bcd_in1=01000011 bcd_in2=01010000 cout=0 sum=10010011
* bcd_in1=01000011 bcd_in2=01010001 cout=0 sum=10010100
* bcd_in1=01000011 bcd_in2=01010010 cout=0 sum=10010101
* bcd_in1=01000011 bcd_in2=01010011 cout=0 sum=10010110
* bcd_in1=01000011 bcd_in2=01010100 cout=0 sum=10010111
* bcd_in1=01000011 bcd_in2=01010101 cout=0 sum=10011000
* bcd_in1=01000011 bcd_in2=01010110 cout=0 sum=10011001
* bcd_in1=01000011 bcd_in2=01010111 cout=1 sum=00000000
* bcd_in1=01000011 bcd_in2=01011000 cout=1 sum=00000001
* bcd_in1=01000011 bcd_in2=01011001 cout=1 sum=00000010
* bcd_in1=01000011 bcd_in2=01100000 cout=1 sum=00000011
* bcd_in1=01000011 bcd_in2=01100001 cout=1 sum=00000100
* bcd_in1=01000011 bcd_in2=01100010 cout=1 sum=00000101
* bcd_in1=01000011 bcd_in2=01100011 cout=1 sum=00000110
* bcd_in1=01000011 bcd_in2=01100100 cout=1 sum=00000111
* bcd_in1=01000011 bcd_in2=01100101 cout=1 sum=00001000
* bcd_in1=01000011 bcd_in2=01100110 cout=1 sum=00001001
* bcd_in1=01000011 bcd_in2=01100111 cout=1 sum=00010000
* bcd_in1=01000011 bcd_in2=01101000 cout=1 sum=00010001
* bcd_in1=01000011 bcd_in2=01101001 cout=1 sum=00010010
* bcd_in1=01000011 bcd_in2=01110000 cout=1 sum=00010011
* bcd_in1=01000011 bcd_in2=01110001 cout=1 sum=00010100
* bcd_in1=01000011 bcd_in2=01110010 cout=1 sum=00010101
* bcd_in1=01000011 bcd_in2=01110011 cout=1 sum=00010110
* bcd_in1=01000011 bcd_in2=01110100 cout=1 sum=00010111
* bcd_in1=01000011 bcd_in2=01110101 cout=1 sum=00011000
* bcd_in1=01000011 bcd_in2=01110110 cout=1 sum=00011001
* bcd_in1=01000011 bcd_in2=01110111 cout=1 sum=00100000
* bcd_in1=01000011 bcd_in2=01111000 cout=1 sum=00100001
* bcd_in1=01000011 bcd_in2=01111001 cout=1 sum=00100010
* bcd_in1=01000011 bcd_in2=10000000 cout=1 sum=00100011
* bcd_in1=01000011 bcd_in2=10000001 cout=1 sum=00100100
* bcd_in1=01000011 bcd_in2=10000010 cout=1 sum=00100101
* bcd_in1=01000011 bcd_in2=10000011 cout=1 sum=00100110
* bcd_in1=01000011 bcd_in2=10000100 cout=1 sum=00100111
* bcd_in1=01000011 bcd_in2=10000101 cout=1 sum=00101000
* bcd_in1=01000011 bcd_in2=10000110 cout=1 sum=00101001
* bcd_in1=01000011 bcd_in2=10000111 cout=1 sum=00110000
* bcd_in1=01000011 bcd_in2=10001000 cout=1 sum=00110001
* bcd_in1=01000011 bcd_in2=10001001 cout=1 sum=00110010
* bcd_in1=01000011 bcd_in2=10010000 cout=1 sum=00110011
* bcd_in1=01000011 bcd_in2=10010001 cout=1 sum=00110100
* bcd_in1=01000011 bcd_in2=10010010 cout=1 sum=00110101
* bcd_in1=01000011 bcd_in2=10010011 cout=1 sum=00110110
* bcd_in1=01000011 bcd_in2=10010100 cout=1 sum=00110111
* bcd_in1=01000011 bcd_in2=10010101 cout=1 sum=00111000
* bcd_in1=01000011 bcd_in2=10010110 cout=1 sum=00111001
* bcd_in1=01000011 bcd_in2=10010111 cout=1 sum=01000000
* bcd_in1=01000011 bcd_in2=10011000 cout=1 sum=01000001
* bcd_in1=01000011 bcd_in2=10011001 cout=1 sum=01000010
* bcd_in1=01000100 bcd_in2=00000000 cout=0 sum=01000100
* bcd_in1=01000100 bcd_in2=00000001 cout=0 sum=01000101
* bcd_in1=01000100 bcd_in2=00000010 cout=0 sum=01000110
* bcd_in1=01000100 bcd_in2=00000011 cout=0 sum=01000111
* bcd_in1=01000100 bcd_in2=00000100 cout=0 sum=01001000
* bcd_in1=01000100 bcd_in2=00000101 cout=0 sum=01001001
* bcd_in1=01000100 bcd_in2=00000110 cout=0 sum=01010000
* bcd_in1=01000100 bcd_in2=00000111 cout=0 sum=01010001
* bcd_in1=01000100 bcd_in2=00001000 cout=0 sum=01010010
* bcd_in1=01000100 bcd_in2=00001001 cout=0 sum=01010011
* bcd_in1=01000100 bcd_in2=00010000 cout=0 sum=01010100
* bcd_in1=01000100 bcd_in2=00010001 cout=0 sum=01010101
* bcd_in1=01000100 bcd_in2=00010010 cout=0 sum=01010110
* bcd_in1=01000100 bcd_in2=00010011 cout=0 sum=01010111
* bcd_in1=01000100 bcd_in2=00010100 cout=0 sum=01011000
* bcd_in1=01000100 bcd_in2=00010101 cout=0 sum=01011001
* bcd_in1=01000100 bcd_in2=00010110 cout=0 sum=01100000
* bcd_in1=01000100 bcd_in2=00010111 cout=0 sum=01100001
* bcd_in1=01000100 bcd_in2=00011000 cout=0 sum=01100010
* bcd_in1=01000100 bcd_in2=00011001 cout=0 sum=01100011
* bcd_in1=01000100 bcd_in2=00100000 cout=0 sum=01100100
* bcd_in1=01000100 bcd_in2=00100001 cout=0 sum=01100101
* bcd_in1=01000100 bcd_in2=00100010 cout=0 sum=01100110
* bcd_in1=01000100 bcd_in2=00100011 cout=0 sum=01100111
* bcd_in1=01000100 bcd_in2=00100100 cout=0 sum=01101000
* bcd_in1=01000100 bcd_in2=00100101 cout=0 sum=01101001
* bcd_in1=01000100 bcd_in2=00100110 cout=0 sum=01110000
* bcd_in1=01000100 bcd_in2=00100111 cout=0 sum=01110001
* bcd_in1=01000100 bcd_in2=00101000 cout=0 sum=01110010
* bcd_in1=01000100 bcd_in2=00101001 cout=0 sum=01110011
* bcd_in1=01000100 bcd_in2=00110000 cout=0 sum=01110100
* bcd_in1=01000100 bcd_in2=00110001 cout=0 sum=01110101
* bcd_in1=01000100 bcd_in2=00110010 cout=0 sum=01110110
* bcd_in1=01000100 bcd_in2=00110011 cout=0 sum=01110111
* bcd_in1=01000100 bcd_in2=00110100 cout=0 sum=01111000
* bcd_in1=01000100 bcd_in2=00110101 cout=0 sum=01111001
* bcd_in1=01000100 bcd_in2=00110110 cout=0 sum=10000000
* bcd_in1=01000100 bcd_in2=00110111 cout=0 sum=10000001
* bcd_in1=01000100 bcd_in2=00111000 cout=0 sum=10000010
* bcd_in1=01000100 bcd_in2=00111001 cout=0 sum=10000011
* bcd_in1=01000100 bcd_in2=01000000 cout=0 sum=10000100
* bcd_in1=01000100 bcd_in2=01000001 cout=0 sum=10000101
* bcd_in1=01000100 bcd_in2=01000010 cout=0 sum=10000110
* bcd_in1=01000100 bcd_in2=01000011 cout=0 sum=10000111
* bcd_in1=01000100 bcd_in2=01000100 cout=0 sum=10001000
* bcd_in1=01000100 bcd_in2=01000101 cout=0 sum=10001001
* bcd_in1=01000100 bcd_in2=01000110 cout=0 sum=10010000
* bcd_in1=01000100 bcd_in2=01000111 cout=0 sum=10010001
* bcd_in1=01000100 bcd_in2=01001000 cout=0 sum=10010010
* bcd_in1=01000100 bcd_in2=01001001 cout=0 sum=10010011
* bcd_in1=01000100 bcd_in2=01010000 cout=0 sum=10010100
* bcd_in1=01000100 bcd_in2=01010001 cout=0 sum=10010101
* bcd_in1=01000100 bcd_in2=01010010 cout=0 sum=10010110
* bcd_in1=01000100 bcd_in2=01010011 cout=0 sum=10010111
* bcd_in1=01000100 bcd_in2=01010100 cout=0 sum=10011000
* bcd_in1=01000100 bcd_in2=01010101 cout=0 sum=10011001
* bcd_in1=01000100 bcd_in2=01010110 cout=1 sum=00000000
* bcd_in1=01000100 bcd_in2=01010111 cout=1 sum=00000001
* bcd_in1=01000100 bcd_in2=01011000 cout=1 sum=00000010
* bcd_in1=01000100 bcd_in2=01011001 cout=1 sum=00000011
* bcd_in1=01000100 bcd_in2=01100000 cout=1 sum=00000100
* bcd_in1=01000100 bcd_in2=01100001 cout=1 sum=00000101
* bcd_in1=01000100 bcd_in2=01100010 cout=1 sum=00000110
* bcd_in1=01000100 bcd_in2=01100011 cout=1 sum=00000111
* bcd_in1=01000100 bcd_in2=01100100 cout=1 sum=00001000
* bcd_in1=01000100 bcd_in2=01100101 cout=1 sum=00001001
* bcd_in1=01000100 bcd_in2=01100110 cout=1 sum=00010000
* bcd_in1=01000100 bcd_in2=01100111 cout=1 sum=00010001
* bcd_in1=01000100 bcd_in2=01101000 cout=1 sum=00010010
* bcd_in1=01000100 bcd_in2=01101001 cout=1 sum=00010011
* bcd_in1=01000100 bcd_in2=01110000 cout=1 sum=00010100
* bcd_in1=01000100 bcd_in2=01110001 cout=1 sum=00010101
* bcd_in1=01000100 bcd_in2=01110010 cout=1 sum=00010110
* bcd_in1=01000100 bcd_in2=01110011 cout=1 sum=00010111
* bcd_in1=01000100 bcd_in2=01110100 cout=1 sum=00011000
* bcd_in1=01000100 bcd_in2=01110101 cout=1 sum=00011001
* bcd_in1=01000100 bcd_in2=01110110 cout=1 sum=00100000
* bcd_in1=01000100 bcd_in2=01110111 cout=1 sum=00100001
* bcd_in1=01000100 bcd_in2=01111000 cout=1 sum=00100010
* bcd_in1=01000100 bcd_in2=01111001 cout=1 sum=00100011
* bcd_in1=01000100 bcd_in2=10000000 cout=1 sum=00100100
* bcd_in1=01000100 bcd_in2=10000001 cout=1 sum=00100101
* bcd_in1=01000100 bcd_in2=10000010 cout=1 sum=00100110
* bcd_in1=01000100 bcd_in2=10000011 cout=1 sum=00100111
* bcd_in1=01000100 bcd_in2=10000100 cout=1 sum=00101000
* bcd_in1=01000100 bcd_in2=10000101 cout=1 sum=00101001
* bcd_in1=01000100 bcd_in2=10000110 cout=1 sum=00110000
* bcd_in1=01000100 bcd_in2=10000111 cout=1 sum=00110001
* bcd_in1=01000100 bcd_in2=10001000 cout=1 sum=00110010
* bcd_in1=01000100 bcd_in2=10001001 cout=1 sum=00110011
* bcd_in1=01000100 bcd_in2=10010000 cout=1 sum=00110100
* bcd_in1=01000100 bcd_in2=10010001 cout=1 sum=00110101
* bcd_in1=01000100 bcd_in2=10010010 cout=1 sum=00110110
* bcd_in1=01000100 bcd_in2=10010011 cout=1 sum=00110111
* bcd_in1=01000100 bcd_in2=10010100 cout=1 sum=00111000
* bcd_in1=01000100 bcd_in2=10010101 cout=1 sum=00111001
* bcd_in1=01000100 bcd_in2=10010110 cout=1 sum=01000000
* bcd_in1=01000100 bcd_in2=10010111 cout=1 sum=01000001
* bcd_in1=01000100 bcd_in2=10011000 cout=1 sum=01000010
* bcd_in1=01000100 bcd_in2=10011001 cout=1 sum=01000011
* bcd_in1=01000101 bcd_in2=00000000 cout=0 sum=01000101
* bcd_in1=01000101 bcd_in2=00000001 cout=0 sum=01000110
* bcd_in1=01000101 bcd_in2=00000010 cout=0 sum=01000111
* bcd_in1=01000101 bcd_in2=00000011 cout=0 sum=01001000
* bcd_in1=01000101 bcd_in2=00000100 cout=0 sum=01001001
* bcd_in1=01000101 bcd_in2=00000101 cout=0 sum=01010000
* bcd_in1=01000101 bcd_in2=00000110 cout=0 sum=01010001
* bcd_in1=01000101 bcd_in2=00000111 cout=0 sum=01010010
* bcd_in1=01000101 bcd_in2=00001000 cout=0 sum=01010011
* bcd_in1=01000101 bcd_in2=00001001 cout=0 sum=01010100
* bcd_in1=01000101 bcd_in2=00010000 cout=0 sum=01010101
* bcd_in1=01000101 bcd_in2=00010001 cout=0 sum=01010110
* bcd_in1=01000101 bcd_in2=00010010 cout=0 sum=01010111
* bcd_in1=01000101 bcd_in2=00010011 cout=0 sum=01011000
* bcd_in1=01000101 bcd_in2=00010100 cout=0 sum=01011001
* bcd_in1=01000101 bcd_in2=00010101 cout=0 sum=01100000
* bcd_in1=01000101 bcd_in2=00010110 cout=0 sum=01100001
* bcd_in1=01000101 bcd_in2=00010111 cout=0 sum=01100010
* bcd_in1=01000101 bcd_in2=00011000 cout=0 sum=01100011
* bcd_in1=01000101 bcd_in2=00011001 cout=0 sum=01100100
* bcd_in1=01000101 bcd_in2=00100000 cout=0 sum=01100101
* bcd_in1=01000101 bcd_in2=00100001 cout=0 sum=01100110
* bcd_in1=01000101 bcd_in2=00100010 cout=0 sum=01100111
* bcd_in1=01000101 bcd_in2=00100011 cout=0 sum=01101000
* bcd_in1=01000101 bcd_in2=00100100 cout=0 sum=01101001
* bcd_in1=01000101 bcd_in2=00100101 cout=0 sum=01110000
* bcd_in1=01000101 bcd_in2=00100110 cout=0 sum=01110001
* bcd_in1=01000101 bcd_in2=00100111 cout=0 sum=01110010
* bcd_in1=01000101 bcd_in2=00101000 cout=0 sum=01110011
* bcd_in1=01000101 bcd_in2=00101001 cout=0 sum=01110100
* bcd_in1=01000101 bcd_in2=00110000 cout=0 sum=01110101
* bcd_in1=01000101 bcd_in2=00110001 cout=0 sum=01110110
* bcd_in1=01000101 bcd_in2=00110010 cout=0 sum=01110111
* bcd_in1=01000101 bcd_in2=00110011 cout=0 sum=01111000
* bcd_in1=01000101 bcd_in2=00110100 cout=0 sum=01111001
* bcd_in1=01000101 bcd_in2=00110101 cout=0 sum=10000000
* bcd_in1=01000101 bcd_in2=00110110 cout=0 sum=10000001
* bcd_in1=01000101 bcd_in2=00110111 cout=0 sum=10000010
* bcd_in1=01000101 bcd_in2=00111000 cout=0 sum=10000011
* bcd_in1=01000101 bcd_in2=00111001 cout=0 sum=10000100
* bcd_in1=01000101 bcd_in2=01000000 cout=0 sum=10000101
* bcd_in1=01000101 bcd_in2=01000001 cout=0 sum=10000110
* bcd_in1=01000101 bcd_in2=01000010 cout=0 sum=10000111
* bcd_in1=01000101 bcd_in2=01000011 cout=0 sum=10001000
* bcd_in1=01000101 bcd_in2=01000100 cout=0 sum=10001001
* bcd_in1=01000101 bcd_in2=01000101 cout=0 sum=10010000
* bcd_in1=01000101 bcd_in2=01000110 cout=0 sum=10010001
* bcd_in1=01000101 bcd_in2=01000111 cout=0 sum=10010010
* bcd_in1=01000101 bcd_in2=01001000 cout=0 sum=10010011
* bcd_in1=01000101 bcd_in2=01001001 cout=0 sum=10010100
* bcd_in1=01000101 bcd_in2=01010000 cout=0 sum=10010101
* bcd_in1=01000101 bcd_in2=01010001 cout=0 sum=10010110
* bcd_in1=01000101 bcd_in2=01010010 cout=0 sum=10010111
* bcd_in1=01000101 bcd_in2=01010011 cout=0 sum=10011000
* bcd_in1=01000101 bcd_in2=01010100 cout=0 sum=10011001
* bcd_in1=01000101 bcd_in2=01010101 cout=1 sum=00000000
* bcd_in1=01000101 bcd_in2=01010110 cout=1 sum=00000001
* bcd_in1=01000101 bcd_in2=01010111 cout=1 sum=00000010
* bcd_in1=01000101 bcd_in2=01011000 cout=1 sum=00000011
* bcd_in1=01000101 bcd_in2=01011001 cout=1 sum=00000100
* bcd_in1=01000101 bcd_in2=01100000 cout=1 sum=00000101
* bcd_in1=01000101 bcd_in2=01100001 cout=1 sum=00000110
* bcd_in1=01000101 bcd_in2=01100010 cout=1 sum=00000111
* bcd_in1=01000101 bcd_in2=01100011 cout=1 sum=00001000
* bcd_in1=01000101 bcd_in2=01100100 cout=1 sum=00001001
* bcd_in1=01000101 bcd_in2=01100101 cout=1 sum=00010000
* bcd_in1=01000101 bcd_in2=01100110 cout=1 sum=00010001
* bcd_in1=01000101 bcd_in2=01100111 cout=1 sum=00010010
* bcd_in1=01000101 bcd_in2=01101000 cout=1 sum=00010011
* bcd_in1=01000101 bcd_in2=01101001 cout=1 sum=00010100
* bcd_in1=01000101 bcd_in2=01110000 cout=1 sum=00010101
* bcd_in1=01000101 bcd_in2=01110001 cout=1 sum=00010110
* bcd_in1=01000101 bcd_in2=01110010 cout=1 sum=00010111
* bcd_in1=01000101 bcd_in2=01110011 cout=1 sum=00011000
* bcd_in1=01000101 bcd_in2=01110100 cout=1 sum=00011001
* bcd_in1=01000101 bcd_in2=01110101 cout=1 sum=00100000
* bcd_in1=01000101 bcd_in2=01110110 cout=1 sum=00100001
* bcd_in1=01000101 bcd_in2=01110111 cout=1 sum=00100010
* bcd_in1=01000101 bcd_in2=01111000 cout=1 sum=00100011
* bcd_in1=01000101 bcd_in2=01111001 cout=1 sum=00100100
* bcd_in1=01000101 bcd_in2=10000000 cout=1 sum=00100101
* bcd_in1=01000101 bcd_in2=10000001 cout=1 sum=00100110
* bcd_in1=01000101 bcd_in2=10000010 cout=1 sum=00100111
* bcd_in1=01000101 bcd_in2=10000011 cout=1 sum=00101000
* bcd_in1=01000101 bcd_in2=10000100 cout=1 sum=00101001
* bcd_in1=01000101 bcd_in2=10000101 cout=1 sum=00110000
* bcd_in1=01000101 bcd_in2=10000110 cout=1 sum=00110001
* bcd_in1=01000101 bcd_in2=10000111 cout=1 sum=00110010
* bcd_in1=01000101 bcd_in2=10001000 cout=1 sum=00110011
* bcd_in1=01000101 bcd_in2=10001001 cout=1 sum=00110100
* bcd_in1=01000101 bcd_in2=10010000 cout=1 sum=00110101
* bcd_in1=01000101 bcd_in2=10010001 cout=1 sum=00110110
* bcd_in1=01000101 bcd_in2=10010010 cout=1 sum=00110111
* bcd_in1=01000101 bcd_in2=10010011 cout=1 sum=00111000
* bcd_in1=01000101 bcd_in2=10010100 cout=1 sum=00111001
* bcd_in1=01000101 bcd_in2=10010101 cout=1 sum=01000000
* bcd_in1=01000101 bcd_in2=10010110 cout=1 sum=01000001
* bcd_in1=01000101 bcd_in2=10010111 cout=1 sum=01000010
* bcd_in1=01000101 bcd_in2=10011000 cout=1 sum=01000011
* bcd_in1=01000101 bcd_in2=10011001 cout=1 sum=01000100
* bcd_in1=01000110 bcd_in2=00000000 cout=0 sum=01000110
* bcd_in1=01000110 bcd_in2=00000001 cout=0 sum=01000111
* bcd_in1=01000110 bcd_in2=00000010 cout=0 sum=01001000
* bcd_in1=01000110 bcd_in2=00000011 cout=0 sum=01001001
* bcd_in1=01000110 bcd_in2=00000100 cout=0 sum=01010000
* bcd_in1=01000110 bcd_in2=00000101 cout=0 sum=01010001
* bcd_in1=01000110 bcd_in2=00000110 cout=0 sum=01010010
* bcd_in1=01000110 bcd_in2=00000111 cout=0 sum=01010011
* bcd_in1=01000110 bcd_in2=00001000 cout=0 sum=01010100
* bcd_in1=01000110 bcd_in2=00001001 cout=0 sum=01010101
* bcd_in1=01000110 bcd_in2=00010000 cout=0 sum=01010110
* bcd_in1=01000110 bcd_in2=00010001 cout=0 sum=01010111
* bcd_in1=01000110 bcd_in2=00010010 cout=0 sum=01011000
* bcd_in1=01000110 bcd_in2=00010011 cout=0 sum=01011001
* bcd_in1=01000110 bcd_in2=00010100 cout=0 sum=01100000
* bcd_in1=01000110 bcd_in2=00010101 cout=0 sum=01100001
* bcd_in1=01000110 bcd_in2=00010110 cout=0 sum=01100010
* bcd_in1=01000110 bcd_in2=00010111 cout=0 sum=01100011
* bcd_in1=01000110 bcd_in2=00011000 cout=0 sum=01100100
* bcd_in1=01000110 bcd_in2=00011001 cout=0 sum=01100101
* bcd_in1=01000110 bcd_in2=00100000 cout=0 sum=01100110
* bcd_in1=01000110 bcd_in2=00100001 cout=0 sum=01100111
* bcd_in1=01000110 bcd_in2=00100010 cout=0 sum=01101000
* bcd_in1=01000110 bcd_in2=00100011 cout=0 sum=01101001
* bcd_in1=01000110 bcd_in2=00100100 cout=0 sum=01110000
* bcd_in1=01000110 bcd_in2=00100101 cout=0 sum=01110001
* bcd_in1=01000110 bcd_in2=00100110 cout=0 sum=01110010
* bcd_in1=01000110 bcd_in2=00100111 cout=0 sum=01110011
* bcd_in1=01000110 bcd_in2=00101000 cout=0 sum=01110100
* bcd_in1=01000110 bcd_in2=00101001 cout=0 sum=01110101
* bcd_in1=01000110 bcd_in2=00110000 cout=0 sum=01110110
* bcd_in1=01000110 bcd_in2=00110001 cout=0 sum=01110111
* bcd_in1=01000110 bcd_in2=00110010 cout=0 sum=01111000
* bcd_in1=01000110 bcd_in2=00110011 cout=0 sum=01111001
* bcd_in1=01000110 bcd_in2=00110100 cout=0 sum=10000000
* bcd_in1=01000110 bcd_in2=00110101 cout=0 sum=10000001
* bcd_in1=01000110 bcd_in2=00110110 cout=0 sum=10000010
* bcd_in1=01000110 bcd_in2=00110111 cout=0 sum=10000011
* bcd_in1=01000110 bcd_in2=00111000 cout=0 sum=10000100
* bcd_in1=01000110 bcd_in2=00111001 cout=0 sum=10000101
* bcd_in1=01000110 bcd_in2=01000000 cout=0 sum=10000110
* bcd_in1=01000110 bcd_in2=01000001 cout=0 sum=10000111
* bcd_in1=01000110 bcd_in2=01000010 cout=0 sum=10001000
* bcd_in1=01000110 bcd_in2=01000011 cout=0 sum=10001001
* bcd_in1=01000110 bcd_in2=01000100 cout=0 sum=10010000
* bcd_in1=01000110 bcd_in2=01000101 cout=0 sum=10010001
* bcd_in1=01000110 bcd_in2=01000110 cout=0 sum=10010010
* bcd_in1=01000110 bcd_in2=01000111 cout=0 sum=10010011
* bcd_in1=01000110 bcd_in2=01001000 cout=0 sum=10010100
* bcd_in1=01000110 bcd_in2=01001001 cout=0 sum=10010101
* bcd_in1=01000110 bcd_in2=01010000 cout=0 sum=10010110
* bcd_in1=01000110 bcd_in2=01010001 cout=0 sum=10010111
* bcd_in1=01000110 bcd_in2=01010010 cout=0 sum=10011000
* bcd_in1=01000110 bcd_in2=01010011 cout=0 sum=10011001
* bcd_in1=01000110 bcd_in2=01010100 cout=1 sum=00000000
* bcd_in1=01000110 bcd_in2=01010101 cout=1 sum=00000001
* bcd_in1=01000110 bcd_in2=01010110 cout=1 sum=00000010
* bcd_in1=01000110 bcd_in2=01010111 cout=1 sum=00000011
* bcd_in1=01000110 bcd_in2=01011000 cout=1 sum=00000100
* bcd_in1=01000110 bcd_in2=01011001 cout=1 sum=00000101
* bcd_in1=01000110 bcd_in2=01100000 cout=1 sum=00000110
* bcd_in1=01000110 bcd_in2=01100001 cout=1 sum=00000111
* bcd_in1=01000110 bcd_in2=01100010 cout=1 sum=00001000
* bcd_in1=01000110 bcd_in2=01100011 cout=1 sum=00001001
* bcd_in1=01000110 bcd_in2=01100100 cout=1 sum=00010000
* bcd_in1=01000110 bcd_in2=01100101 cout=1 sum=00010001
* bcd_in1=01000110 bcd_in2=01100110 cout=1 sum=00010010
* bcd_in1=01000110 bcd_in2=01100111 cout=1 sum=00010011
* bcd_in1=01000110 bcd_in2=01101000 cout=1 sum=00010100
* bcd_in1=01000110 bcd_in2=01101001 cout=1 sum=00010101
* bcd_in1=01000110 bcd_in2=01110000 cout=1 sum=00010110
* bcd_in1=01000110 bcd_in2=01110001 cout=1 sum=00010111
* bcd_in1=01000110 bcd_in2=01110010 cout=1 sum=00011000
* bcd_in1=01000110 bcd_in2=01110011 cout=1 sum=00011001
* bcd_in1=01000110 bcd_in2=01110100 cout=1 sum=00100000
* bcd_in1=01000110 bcd_in2=01110101 cout=1 sum=00100001
* bcd_in1=01000110 bcd_in2=01110110 cout=1 sum=00100010
* bcd_in1=01000110 bcd_in2=01110111 cout=1 sum=00100011
* bcd_in1=01000110 bcd_in2=01111000 cout=1 sum=00100100
* bcd_in1=01000110 bcd_in2=01111001 cout=1 sum=00100101
* bcd_in1=01000110 bcd_in2=10000000 cout=1 sum=00100110
* bcd_in1=01000110 bcd_in2=10000001 cout=1 sum=00100111
* bcd_in1=01000110 bcd_in2=10000010 cout=1 sum=00101000
* bcd_in1=01000110 bcd_in2=10000011 cout=1 sum=00101001
* bcd_in1=01000110 bcd_in2=10000100 cout=1 sum=00110000
* bcd_in1=01000110 bcd_in2=10000101 cout=1 sum=00110001
* bcd_in1=01000110 bcd_in2=10000110 cout=1 sum=00110010
* bcd_in1=01000110 bcd_in2=10000111 cout=1 sum=00110011
* bcd_in1=01000110 bcd_in2=10001000 cout=1 sum=00110100
* bcd_in1=01000110 bcd_in2=10001001 cout=1 sum=00110101
* bcd_in1=01000110 bcd_in2=10010000 cout=1 sum=00110110
* bcd_in1=01000110 bcd_in2=10010001 cout=1 sum=00110111
* bcd_in1=01000110 bcd_in2=10010010 cout=1 sum=00111000
* bcd_in1=01000110 bcd_in2=10010011 cout=1 sum=00111001
* bcd_in1=01000110 bcd_in2=10010100 cout=1 sum=01000000
* bcd_in1=01000110 bcd_in2=10010101 cout=1 sum=01000001
* bcd_in1=01000110 bcd_in2=10010110 cout=1 sum=01000010
* bcd_in1=01000110 bcd_in2=10010111 cout=1 sum=01000011
* bcd_in1=01000110 bcd_in2=10011000 cout=1 sum=01000100
* bcd_in1=01000110 bcd_in2=10011001 cout=1 sum=01000101
* bcd_in1=01000111 bcd_in2=00000000 cout=0 sum=01000111
* bcd_in1=01000111 bcd_in2=00000001 cout=0 sum=01001000
* bcd_in1=01000111 bcd_in2=00000010 cout=0 sum=01001001
* bcd_in1=01000111 bcd_in2=00000011 cout=0 sum=01010000
* bcd_in1=01000111 bcd_in2=00000100 cout=0 sum=01010001
* bcd_in1=01000111 bcd_in2=00000101 cout=0 sum=01010010
* bcd_in1=01000111 bcd_in2=00000110 cout=0 sum=01010011
* bcd_in1=01000111 bcd_in2=00000111 cout=0 sum=01010100
* bcd_in1=01000111 bcd_in2=00001000 cout=0 sum=01010101
* bcd_in1=01000111 bcd_in2=00001001 cout=0 sum=01010110
* bcd_in1=01000111 bcd_in2=00010000 cout=0 sum=01010111
* bcd_in1=01000111 bcd_in2=00010001 cout=0 sum=01011000
* bcd_in1=01000111 bcd_in2=00010010 cout=0 sum=01011001
* bcd_in1=01000111 bcd_in2=00010011 cout=0 sum=01100000
* bcd_in1=01000111 bcd_in2=00010100 cout=0 sum=01100001
* bcd_in1=01000111 bcd_in2=00010101 cout=0 sum=01100010
* bcd_in1=01000111 bcd_in2=00010110 cout=0 sum=01100011
* bcd_in1=01000111 bcd_in2=00010111 cout=0 sum=01100100
* bcd_in1=01000111 bcd_in2=00011000 cout=0 sum=01100101
* bcd_in1=01000111 bcd_in2=00011001 cout=0 sum=01100110
* bcd_in1=01000111 bcd_in2=00100000 cout=0 sum=01100111
* bcd_in1=01000111 bcd_in2=00100001 cout=0 sum=01101000
* bcd_in1=01000111 bcd_in2=00100010 cout=0 sum=01101001
* bcd_in1=01000111 bcd_in2=00100011 cout=0 sum=01110000
* bcd_in1=01000111 bcd_in2=00100100 cout=0 sum=01110001
* bcd_in1=01000111 bcd_in2=00100101 cout=0 sum=01110010
* bcd_in1=01000111 bcd_in2=00100110 cout=0 sum=01110011
* bcd_in1=01000111 bcd_in2=00100111 cout=0 sum=01110100
* bcd_in1=01000111 bcd_in2=00101000 cout=0 sum=01110101
* bcd_in1=01000111 bcd_in2=00101001 cout=0 sum=01110110
* bcd_in1=01000111 bcd_in2=00110000 cout=0 sum=01110111
* bcd_in1=01000111 bcd_in2=00110001 cout=0 sum=01111000
* bcd_in1=01000111 bcd_in2=00110010 cout=0 sum=01111001
* bcd_in1=01000111 bcd_in2=00110011 cout=0 sum=10000000
* bcd_in1=01000111 bcd_in2=00110100 cout=0 sum=10000001
* bcd_in1=01000111 bcd_in2=00110101 cout=0 sum=10000010
* bcd_in1=01000111 bcd_in2=00110110 cout=0 sum=10000011
* bcd_in1=01000111 bcd_in2=00110111 cout=0 sum=10000100
* bcd_in1=01000111 bcd_in2=00111000 cout=0 sum=10000101
* bcd_in1=01000111 bcd_in2=00111001 cout=0 sum=10000110
* bcd_in1=01000111 bcd_in2=01000000 cout=0 sum=10000111
* bcd_in1=01000111 bcd_in2=01000001 cout=0 sum=10001000
* bcd_in1=01000111 bcd_in2=01000010 cout=0 sum=10001001
* bcd_in1=01000111 bcd_in2=01000011 cout=0 sum=10010000
* bcd_in1=01000111 bcd_in2=01000100 cout=0 sum=10010001
* bcd_in1=01000111 bcd_in2=01000101 cout=0 sum=10010010
* bcd_in1=01000111 bcd_in2=01000110 cout=0 sum=10010011
* bcd_in1=01000111 bcd_in2=01000111 cout=0 sum=10010100
* bcd_in1=01000111 bcd_in2=01001000 cout=0 sum=10010101
* bcd_in1=01000111 bcd_in2=01001001 cout=0 sum=10010110
* bcd_in1=01000111 bcd_in2=01010000 cout=0 sum=10010111
* bcd_in1=01000111 bcd_in2=01010001 cout=0 sum=10011000
* bcd_in1=01000111 bcd_in2=01010010 cout=0 sum=10011001
* bcd_in1=01000111 bcd_in2=01010011 cout=1 sum=00000000
* bcd_in1=01000111 bcd_in2=01010100 cout=1 sum=00000001
* bcd_in1=01000111 bcd_in2=01010101 cout=1 sum=00000010
* bcd_in1=01000111 bcd_in2=01010110 cout=1 sum=00000011
* bcd_in1=01000111 bcd_in2=01010111 cout=1 sum=00000100
* bcd_in1=01000111 bcd_in2=01011000 cout=1 sum=00000101
* bcd_in1=01000111 bcd_in2=01011001 cout=1 sum=00000110
* bcd_in1=01000111 bcd_in2=01100000 cout=1 sum=00000111
* bcd_in1=01000111 bcd_in2=01100001 cout=1 sum=00001000
* bcd_in1=01000111 bcd_in2=01100010 cout=1 sum=00001001
* bcd_in1=01000111 bcd_in2=01100011 cout=1 sum=00010000
* bcd_in1=01000111 bcd_in2=01100100 cout=1 sum=00010001
* bcd_in1=01000111 bcd_in2=01100101 cout=1 sum=00010010
* bcd_in1=01000111 bcd_in2=01100110 cout=1 sum=00010011
* bcd_in1=01000111 bcd_in2=01100111 cout=1 sum=00010100
* bcd_in1=01000111 bcd_in2=01101000 cout=1 sum=00010101
* bcd_in1=01000111 bcd_in2=01101001 cout=1 sum=00010110
* bcd_in1=01000111 bcd_in2=01110000 cout=1 sum=00010111
* bcd_in1=01000111 bcd_in2=01110001 cout=1 sum=00011000
* bcd_in1=01000111 bcd_in2=01110010 cout=1 sum=00011001
* bcd_in1=01000111 bcd_in2=01110011 cout=1 sum=00100000
* bcd_in1=01000111 bcd_in2=01110100 cout=1 sum=00100001
* bcd_in1=01000111 bcd_in2=01110101 cout=1 sum=00100010
* bcd_in1=01000111 bcd_in2=01110110 cout=1 sum=00100011
* bcd_in1=01000111 bcd_in2=01110111 cout=1 sum=00100100
* bcd_in1=01000111 bcd_in2=01111000 cout=1 sum=00100101
* bcd_in1=01000111 bcd_in2=01111001 cout=1 sum=00100110
* bcd_in1=01000111 bcd_in2=10000000 cout=1 sum=00100111
* bcd_in1=01000111 bcd_in2=10000001 cout=1 sum=00101000
* bcd_in1=01000111 bcd_in2=10000010 cout=1 sum=00101001
* bcd_in1=01000111 bcd_in2=10000011 cout=1 sum=00110000
* bcd_in1=01000111 bcd_in2=10000100 cout=1 sum=00110001
* bcd_in1=01000111 bcd_in2=10000101 cout=1 sum=00110010
* bcd_in1=01000111 bcd_in2=10000110 cout=1 sum=00110011
* bcd_in1=01000111 bcd_in2=10000111 cout=1 sum=00110100
* bcd_in1=01000111 bcd_in2=10001000 cout=1 sum=00110101
* bcd_in1=01000111 bcd_in2=10001001 cout=1 sum=00110110
* bcd_in1=01000111 bcd_in2=10010000 cout=1 sum=00110111
* bcd_in1=01000111 bcd_in2=10010001 cout=1 sum=00111000
* bcd_in1=01000111 bcd_in2=10010010 cout=1 sum=00111001
* bcd_in1=01000111 bcd_in2=10010011 cout=1 sum=01000000
* bcd_in1=01000111 bcd_in2=10010100 cout=1 sum=01000001
* bcd_in1=01000111 bcd_in2=10010101 cout=1 sum=01000010
* bcd_in1=01000111 bcd_in2=10010110 cout=1 sum=01000011
* bcd_in1=01000111 bcd_in2=10010111 cout=1 sum=01000100
* bcd_in1=01000111 bcd_in2=10011000 cout=1 sum=01000101
* bcd_in1=01000111 bcd_in2=10011001 cout=1 sum=01000110
* bcd_in1=01001000 bcd_in2=00000000 cout=0 sum=01001000
* bcd_in1=01001000 bcd_in2=00000001 cout=0 sum=01001001
* bcd_in1=01001000 bcd_in2=00000010 cout=0 sum=01010000
* bcd_in1=01001000 bcd_in2=00000011 cout=0 sum=01010001
* bcd_in1=01001000 bcd_in2=00000100 cout=0 sum=01010010
* bcd_in1=01001000 bcd_in2=00000101 cout=0 sum=01010011
* bcd_in1=01001000 bcd_in2=00000110 cout=0 sum=01010100
* bcd_in1=01001000 bcd_in2=00000111 cout=0 sum=01010101
* bcd_in1=01001000 bcd_in2=00001000 cout=0 sum=01010110
* bcd_in1=01001000 bcd_in2=00001001 cout=0 sum=01010111
* bcd_in1=01001000 bcd_in2=00010000 cout=0 sum=01011000
* bcd_in1=01001000 bcd_in2=00010001 cout=0 sum=01011001
* bcd_in1=01001000 bcd_in2=00010010 cout=0 sum=01100000
* bcd_in1=01001000 bcd_in2=00010011 cout=0 sum=01100001
* bcd_in1=01001000 bcd_in2=00010100 cout=0 sum=01100010
* bcd_in1=01001000 bcd_in2=00010101 cout=0 sum=01100011
* bcd_in1=01001000 bcd_in2=00010110 cout=0 sum=01100100
* bcd_in1=01001000 bcd_in2=00010111 cout=0 sum=01100101
* bcd_in1=01001000 bcd_in2=00011000 cout=0 sum=01100110
* bcd_in1=01001000 bcd_in2=00011001 cout=0 sum=01100111
* bcd_in1=01001000 bcd_in2=00100000 cout=0 sum=01101000
* bcd_in1=01001000 bcd_in2=00100001 cout=0 sum=01101001
* bcd_in1=01001000 bcd_in2=00100010 cout=0 sum=01110000
* bcd_in1=01001000 bcd_in2=00100011 cout=0 sum=01110001
* bcd_in1=01001000 bcd_in2=00100100 cout=0 sum=01110010
* bcd_in1=01001000 bcd_in2=00100101 cout=0 sum=01110011
* bcd_in1=01001000 bcd_in2=00100110 cout=0 sum=01110100
* bcd_in1=01001000 bcd_in2=00100111 cout=0 sum=01110101
* bcd_in1=01001000 bcd_in2=00101000 cout=0 sum=01110110
* bcd_in1=01001000 bcd_in2=00101001 cout=0 sum=01110111
* bcd_in1=01001000 bcd_in2=00110000 cout=0 sum=01111000
* bcd_in1=01001000 bcd_in2=00110001 cout=0 sum=01111001
* bcd_in1=01001000 bcd_in2=00110010 cout=0 sum=10000000
* bcd_in1=01001000 bcd_in2=00110011 cout=0 sum=10000001
* bcd_in1=01001000 bcd_in2=00110100 cout=0 sum=10000010
* bcd_in1=01001000 bcd_in2=00110101 cout=0 sum=10000011
* bcd_in1=01001000 bcd_in2=00110110 cout=0 sum=10000100
* bcd_in1=01001000 bcd_in2=00110111 cout=0 sum=10000101
* bcd_in1=01001000 bcd_in2=00111000 cout=0 sum=10000110
* bcd_in1=01001000 bcd_in2=00111001 cout=0 sum=10000111
* bcd_in1=01001000 bcd_in2=01000000 cout=0 sum=10001000
* bcd_in1=01001000 bcd_in2=01000001 cout=0 sum=10001001
* bcd_in1=01001000 bcd_in2=01000010 cout=0 sum=10010000
* bcd_in1=01001000 bcd_in2=01000011 cout=0 sum=10010001
* bcd_in1=01001000 bcd_in2=01000100 cout=0 sum=10010010
* bcd_in1=01001000 bcd_in2=01000101 cout=0 sum=10010011
* bcd_in1=01001000 bcd_in2=01000110 cout=0 sum=10010100
* bcd_in1=01001000 bcd_in2=01000111 cout=0 sum=10010101
* bcd_in1=01001000 bcd_in2=01001000 cout=0 sum=10010110
* bcd_in1=01001000 bcd_in2=01001001 cout=0 sum=10010111
* bcd_in1=01001000 bcd_in2=01010000 cout=0 sum=10011000
* bcd_in1=01001000 bcd_in2=01010001 cout=0 sum=10011001
* bcd_in1=01001000 bcd_in2=01010010 cout=1 sum=00000000
* bcd_in1=01001000 bcd_in2=01010011 cout=1 sum=00000001
* bcd_in1=01001000 bcd_in2=01010100 cout=1 sum=00000010
* bcd_in1=01001000 bcd_in2=01010101 cout=1 sum=00000011
* bcd_in1=01001000 bcd_in2=01010110 cout=1 sum=00000100
* bcd_in1=01001000 bcd_in2=01010111 cout=1 sum=00000101
* bcd_in1=01001000 bcd_in2=01011000 cout=1 sum=00000110
* bcd_in1=01001000 bcd_in2=01011001 cout=1 sum=00000111
* bcd_in1=01001000 bcd_in2=01100000 cout=1 sum=00001000
* bcd_in1=01001000 bcd_in2=01100001 cout=1 sum=00001001
* bcd_in1=01001000 bcd_in2=01100010 cout=1 sum=00010000
* bcd_in1=01001000 bcd_in2=01100011 cout=1 sum=00010001
* bcd_in1=01001000 bcd_in2=01100100 cout=1 sum=00010010
* bcd_in1=01001000 bcd_in2=01100101 cout=1 sum=00010011
* bcd_in1=01001000 bcd_in2=01100110 cout=1 sum=00010100
* bcd_in1=01001000 bcd_in2=01100111 cout=1 sum=00010101
* bcd_in1=01001000 bcd_in2=01101000 cout=1 sum=00010110
* bcd_in1=01001000 bcd_in2=01101001 cout=1 sum=00010111
* bcd_in1=01001000 bcd_in2=01110000 cout=1 sum=00011000
* bcd_in1=01001000 bcd_in2=01110001 cout=1 sum=00011001
* bcd_in1=01001000 bcd_in2=01110010 cout=1 sum=00100000
* bcd_in1=01001000 bcd_in2=01110011 cout=1 sum=00100001
* bcd_in1=01001000 bcd_in2=01110100 cout=1 sum=00100010
* bcd_in1=01001000 bcd_in2=01110101 cout=1 sum=00100011
* bcd_in1=01001000 bcd_in2=01110110 cout=1 sum=00100100
* bcd_in1=01001000 bcd_in2=01110111 cout=1 sum=00100101
* bcd_in1=01001000 bcd_in2=01111000 cout=1 sum=00100110
* bcd_in1=01001000 bcd_in2=01111001 cout=1 sum=00100111
* bcd_in1=01001000 bcd_in2=10000000 cout=1 sum=00101000
* bcd_in1=01001000 bcd_in2=10000001 cout=1 sum=00101001
* bcd_in1=01001000 bcd_in2=10000010 cout=1 sum=00110000
* bcd_in1=01001000 bcd_in2=10000011 cout=1 sum=00110001
* bcd_in1=01001000 bcd_in2=10000100 cout=1 sum=00110010
* bcd_in1=01001000 bcd_in2=10000101 cout=1 sum=00110011
* bcd_in1=01001000 bcd_in2=10000110 cout=1 sum=00110100
* bcd_in1=01001000 bcd_in2=10000111 cout=1 sum=00110101
* bcd_in1=01001000 bcd_in2=10001000 cout=1 sum=00110110
* bcd_in1=01001000 bcd_in2=10001001 cout=1 sum=00110111
* bcd_in1=01001000 bcd_in2=10010000 cout=1 sum=00111000
* bcd_in1=01001000 bcd_in2=10010001 cout=1 sum=00111001
* bcd_in1=01001000 bcd_in2=10010010 cout=1 sum=01000000
* bcd_in1=01001000 bcd_in2=10010011 cout=1 sum=01000001
* bcd_in1=01001000 bcd_in2=10010100 cout=1 sum=01000010
* bcd_in1=01001000 bcd_in2=10010101 cout=1 sum=01000011
* bcd_in1=01001000 bcd_in2=10010110 cout=1 sum=01000100
* bcd_in1=01001000 bcd_in2=10010111 cout=1 sum=01000101
* bcd_in1=01001000 bcd_in2=10011000 cout=1 sum=01000110
* bcd_in1=01001000 bcd_in2=10011001 cout=1 sum=01000111
* bcd_in1=01001001 bcd_in2=00000000 cout=0 sum=01001001
* bcd_in1=01001001 bcd_in2=00000001 cout=0 sum=01010000
* bcd_in1=01001001 bcd_in2=00000010 cout=0 sum=01010001
* bcd_in1=01001001 bcd_in2=00000011 cout=0 sum=01010010
* bcd_in1=01001001 bcd_in2=00000100 cout=0 sum=01010011
* bcd_in1=01001001 bcd_in2=00000101 cout=0 sum=01010100
* bcd_in1=01001001 bcd_in2=00000110 cout=0 sum=01010101
* bcd_in1=01001001 bcd_in2=00000111 cout=0 sum=01010110
* bcd_in1=01001001 bcd_in2=00001000 cout=0 sum=01010111
* bcd_in1=01001001 bcd_in2=00001001 cout=0 sum=01011000
* bcd_in1=01001001 bcd_in2=00010000 cout=0 sum=01011001
* bcd_in1=01001001 bcd_in2=00010001 cout=0 sum=01100000
* bcd_in1=01001001 bcd_in2=00010010 cout=0 sum=01100001
* bcd_in1=01001001 bcd_in2=00010011 cout=0 sum=01100010
* bcd_in1=01001001 bcd_in2=00010100 cout=0 sum=01100011
* bcd_in1=01001001 bcd_in2=00010101 cout=0 sum=01100100
* bcd_in1=01001001 bcd_in2=00010110 cout=0 sum=01100101
* bcd_in1=01001001 bcd_in2=00010111 cout=0 sum=01100110
* bcd_in1=01001001 bcd_in2=00011000 cout=0 sum=01100111
* bcd_in1=01001001 bcd_in2=00011001 cout=0 sum=01101000
* bcd_in1=01001001 bcd_in2=00100000 cout=0 sum=01101001
* bcd_in1=01001001 bcd_in2=00100001 cout=0 sum=01110000
* bcd_in1=01001001 bcd_in2=00100010 cout=0 sum=01110001
* bcd_in1=01001001 bcd_in2=00100011 cout=0 sum=01110010
* bcd_in1=01001001 bcd_in2=00100100 cout=0 sum=01110011
* bcd_in1=01001001 bcd_in2=00100101 cout=0 sum=01110100
* bcd_in1=01001001 bcd_in2=00100110 cout=0 sum=01110101
* bcd_in1=01001001 bcd_in2=00100111 cout=0 sum=01110110
* bcd_in1=01001001 bcd_in2=00101000 cout=0 sum=01110111
* bcd_in1=01001001 bcd_in2=00101001 cout=0 sum=01111000
* bcd_in1=01001001 bcd_in2=00110000 cout=0 sum=01111001
* bcd_in1=01001001 bcd_in2=00110001 cout=0 sum=10000000
* bcd_in1=01001001 bcd_in2=00110010 cout=0 sum=10000001
* bcd_in1=01001001 bcd_in2=00110011 cout=0 sum=10000010
* bcd_in1=01001001 bcd_in2=00110100 cout=0 sum=10000011
* bcd_in1=01001001 bcd_in2=00110101 cout=0 sum=10000100
* bcd_in1=01001001 bcd_in2=00110110 cout=0 sum=10000101
* bcd_in1=01001001 bcd_in2=00110111 cout=0 sum=10000110
* bcd_in1=01001001 bcd_in2=00111000 cout=0 sum=10000111
* bcd_in1=01001001 bcd_in2=00111001 cout=0 sum=10001000
* bcd_in1=01001001 bcd_in2=01000000 cout=0 sum=10001001
* bcd_in1=01001001 bcd_in2=01000001 cout=0 sum=10010000
* bcd_in1=01001001 bcd_in2=01000010 cout=0 sum=10010001
* bcd_in1=01001001 bcd_in2=01000011 cout=0 sum=10010010
* bcd_in1=01001001 bcd_in2=01000100 cout=0 sum=10010011
* bcd_in1=01001001 bcd_in2=01000101 cout=0 sum=10010100
* bcd_in1=01001001 bcd_in2=01000110 cout=0 sum=10010101
* bcd_in1=01001001 bcd_in2=01000111 cout=0 sum=10010110
* bcd_in1=01001001 bcd_in2=01001000 cout=0 sum=10010111
* bcd_in1=01001001 bcd_in2=01001001 cout=0 sum=10011000
* bcd_in1=01001001 bcd_in2=01010000 cout=0 sum=10011001
* bcd_in1=01001001 bcd_in2=01010001 cout=1 sum=00000000
* bcd_in1=01001001 bcd_in2=01010010 cout=1 sum=00000001
* bcd_in1=01001001 bcd_in2=01010011 cout=1 sum=00000010
* bcd_in1=01001001 bcd_in2=01010100 cout=1 sum=00000011
* bcd_in1=01001001 bcd_in2=01010101 cout=1 sum=00000100
* bcd_in1=01001001 bcd_in2=01010110 cout=1 sum=00000101
* bcd_in1=01001001 bcd_in2=01010111 cout=1 sum=00000110
* bcd_in1=01001001 bcd_in2=01011000 cout=1 sum=00000111
* bcd_in1=01001001 bcd_in2=01011001 cout=1 sum=00001000
* bcd_in1=01001001 bcd_in2=01100000 cout=1 sum=00001001
* bcd_in1=01001001 bcd_in2=01100001 cout=1 sum=00010000
* bcd_in1=01001001 bcd_in2=01100010 cout=1 sum=00010001
* bcd_in1=01001001 bcd_in2=01100011 cout=1 sum=00010010
* bcd_in1=01001001 bcd_in2=01100100 cout=1 sum=00010011
* bcd_in1=01001001 bcd_in2=01100101 cout=1 sum=00010100
* bcd_in1=01001001 bcd_in2=01100110 cout=1 sum=00010101
* bcd_in1=01001001 bcd_in2=01100111 cout=1 sum=00010110
* bcd_in1=01001001 bcd_in2=01101000 cout=1 sum=00010111
* bcd_in1=01001001 bcd_in2=01101001 cout=1 sum=00011000
* bcd_in1=01001001 bcd_in2=01110000 cout=1 sum=00011001
* bcd_in1=01001001 bcd_in2=01110001 cout=1 sum=00100000
* bcd_in1=01001001 bcd_in2=01110010 cout=1 sum=00100001
* bcd_in1=01001001 bcd_in2=01110011 cout=1 sum=00100010
* bcd_in1=01001001 bcd_in2=01110100 cout=1 sum=00100011
* bcd_in1=01001001 bcd_in2=01110101 cout=1 sum=00100100
* bcd_in1=01001001 bcd_in2=01110110 cout=1 sum=00100101
* bcd_in1=01001001 bcd_in2=01110111 cout=1 sum=00100110
* bcd_in1=01001001 bcd_in2=01111000 cout=1 sum=00100111
* bcd_in1=01001001 bcd_in2=01111001 cout=1 sum=00101000
* bcd_in1=01001001 bcd_in2=10000000 cout=1 sum=00101001
* bcd_in1=01001001 bcd_in2=10000001 cout=1 sum=00110000
* bcd_in1=01001001 bcd_in2=10000010 cout=1 sum=00110001
* bcd_in1=01001001 bcd_in2=10000011 cout=1 sum=00110010
* bcd_in1=01001001 bcd_in2=10000100 cout=1 sum=00110011
* bcd_in1=01001001 bcd_in2=10000101 cout=1 sum=00110100
* bcd_in1=01001001 bcd_in2=10000110 cout=1 sum=00110101
* bcd_in1=01001001 bcd_in2=10000111 cout=1 sum=00110110
* bcd_in1=01001001 bcd_in2=10001000 cout=1 sum=00110111
* bcd_in1=01001001 bcd_in2=10001001 cout=1 sum=00111000
* bcd_in1=01001001 bcd_in2=10010000 cout=1 sum=00111001
* bcd_in1=01001001 bcd_in2=10010001 cout=1 sum=01000000
* bcd_in1=01001001 bcd_in2=10010010 cout=1 sum=01000001
* bcd_in1=01001001 bcd_in2=10010011 cout=1 sum=01000010
* bcd_in1=01001001 bcd_in2=10010100 cout=1 sum=01000011
* bcd_in1=01001001 bcd_in2=10010101 cout=1 sum=01000100
* bcd_in1=01001001 bcd_in2=10010110 cout=1 sum=01000101
* bcd_in1=01001001 bcd_in2=10010111 cout=1 sum=01000110
* bcd_in1=01001001 bcd_in2=10011000 cout=1 sum=01000111
* bcd_in1=01001001 bcd_in2=10011001 cout=1 sum=01001000
* bcd_in1=01010000 bcd_in2=00000000 cout=0 sum=01010000
* bcd_in1=01010000 bcd_in2=00000001 cout=0 sum=01010001
* bcd_in1=01010000 bcd_in2=00000010 cout=0 sum=01010010
* bcd_in1=01010000 bcd_in2=00000011 cout=0 sum=01010011
* bcd_in1=01010000 bcd_in2=00000100 cout=0 sum=01010100
* bcd_in1=01010000 bcd_in2=00000101 cout=0 sum=01010101
* bcd_in1=01010000 bcd_in2=00000110 cout=0 sum=01010110
* bcd_in1=01010000 bcd_in2=00000111 cout=0 sum=01010111
* bcd_in1=01010000 bcd_in2=00001000 cout=0 sum=01011000
* bcd_in1=01010000 bcd_in2=00001001 cout=0 sum=01011001
* bcd_in1=01010000 bcd_in2=00010000 cout=0 sum=01100000
* bcd_in1=01010000 bcd_in2=00010001 cout=0 sum=01100001
* bcd_in1=01010000 bcd_in2=00010010 cout=0 sum=01100010
* bcd_in1=01010000 bcd_in2=00010011 cout=0 sum=01100011
* bcd_in1=01010000 bcd_in2=00010100 cout=0 sum=01100100
* bcd_in1=01010000 bcd_in2=00010101 cout=0 sum=01100101
* bcd_in1=01010000 bcd_in2=00010110 cout=0 sum=01100110
* bcd_in1=01010000 bcd_in2=00010111 cout=0 sum=01100111
* bcd_in1=01010000 bcd_in2=00011000 cout=0 sum=01101000
* bcd_in1=01010000 bcd_in2=00011001 cout=0 sum=01101001
* bcd_in1=01010000 bcd_in2=00100000 cout=0 sum=01110000
* bcd_in1=01010000 bcd_in2=00100001 cout=0 sum=01110001
* bcd_in1=01010000 bcd_in2=00100010 cout=0 sum=01110010
* bcd_in1=01010000 bcd_in2=00100011 cout=0 sum=01110011
* bcd_in1=01010000 bcd_in2=00100100 cout=0 sum=01110100
* bcd_in1=01010000 bcd_in2=00100101 cout=0 sum=01110101
* bcd_in1=01010000 bcd_in2=00100110 cout=0 sum=01110110
* bcd_in1=01010000 bcd_in2=00100111 cout=0 sum=01110111
* bcd_in1=01010000 bcd_in2=00101000 cout=0 sum=01111000
* bcd_in1=01010000 bcd_in2=00101001 cout=0 sum=01111001
* bcd_in1=01010000 bcd_in2=00110000 cout=0 sum=10000000
* bcd_in1=01010000 bcd_in2=00110001 cout=0 sum=10000001
* bcd_in1=01010000 bcd_in2=00110010 cout=0 sum=10000010
* bcd_in1=01010000 bcd_in2=00110011 cout=0 sum=10000011
* bcd_in1=01010000 bcd_in2=00110100 cout=0 sum=10000100
* bcd_in1=01010000 bcd_in2=00110101 cout=0 sum=10000101
* bcd_in1=01010000 bcd_in2=00110110 cout=0 sum=10000110
* bcd_in1=01010000 bcd_in2=00110111 cout=0 sum=10000111
* bcd_in1=01010000 bcd_in2=00111000 cout=0 sum=10001000
* bcd_in1=01010000 bcd_in2=00111001 cout=0 sum=10001001
* bcd_in1=01010000 bcd_in2=01000000 cout=0 sum=10010000
* bcd_in1=01010000 bcd_in2=01000001 cout=0 sum=10010001
* bcd_in1=01010000 bcd_in2=01000010 cout=0 sum=10010010
* bcd_in1=01010000 bcd_in2=01000011 cout=0 sum=10010011
* bcd_in1=01010000 bcd_in2=01000100 cout=0 sum=10010100
* bcd_in1=01010000 bcd_in2=01000101 cout=0 sum=10010101
* bcd_in1=01010000 bcd_in2=01000110 cout=0 sum=10010110
* bcd_in1=01010000 bcd_in2=01000111 cout=0 sum=10010111
* bcd_in1=01010000 bcd_in2=01001000 cout=0 sum=10011000
* bcd_in1=01010000 bcd_in2=01001001 cout=0 sum=10011001
* bcd_in1=01010000 bcd_in2=01010000 cout=1 sum=00000000
* bcd_in1=01010000 bcd_in2=01010001 cout=1 sum=00000001
* bcd_in1=01010000 bcd_in2=01010010 cout=1 sum=00000010
* bcd_in1=01010000 bcd_in2=01010011 cout=1 sum=00000011
* bcd_in1=01010000 bcd_in2=01010100 cout=1 sum=00000100
* bcd_in1=01010000 bcd_in2=01010101 cout=1 sum=00000101
* bcd_in1=01010000 bcd_in2=01010110 cout=1 sum=00000110
* bcd_in1=01010000 bcd_in2=01010111 cout=1 sum=00000111
* bcd_in1=01010000 bcd_in2=01011000 cout=1 sum=00001000
* bcd_in1=01010000 bcd_in2=01011001 cout=1 sum=00001001
* bcd_in1=01010000 bcd_in2=01100000 cout=1 sum=00010000
* bcd_in1=01010000 bcd_in2=01100001 cout=1 sum=00010001
* bcd_in1=01010000 bcd_in2=01100010 cout=1 sum=00010010
* bcd_in1=01010000 bcd_in2=01100011 cout=1 sum=00010011
* bcd_in1=01010000 bcd_in2=01100100 cout=1 sum=00010100
* bcd_in1=01010000 bcd_in2=01100101 cout=1 sum=00010101
* bcd_in1=01010000 bcd_in2=01100110 cout=1 sum=00010110
* bcd_in1=01010000 bcd_in2=01100111 cout=1 sum=00010111
* bcd_in1=01010000 bcd_in2=01101000 cout=1 sum=00011000
* bcd_in1=01010000 bcd_in2=01101001 cout=1 sum=00011001
* bcd_in1=01010000 bcd_in2=01110000 cout=1 sum=00100000
* bcd_in1=01010000 bcd_in2=01110001 cout=1 sum=00100001
* bcd_in1=01010000 bcd_in2=01110010 cout=1 sum=00100010
* bcd_in1=01010000 bcd_in2=01110011 cout=1 sum=00100011
* bcd_in1=01010000 bcd_in2=01110100 cout=1 sum=00100100
* bcd_in1=01010000 bcd_in2=01110101 cout=1 sum=00100101
* bcd_in1=01010000 bcd_in2=01110110 cout=1 sum=00100110
* bcd_in1=01010000 bcd_in2=01110111 cout=1 sum=00100111
* bcd_in1=01010000 bcd_in2=01111000 cout=1 sum=00101000
* bcd_in1=01010000 bcd_in2=01111001 cout=1 sum=00101001
* bcd_in1=01010000 bcd_in2=10000000 cout=1 sum=00110000
* bcd_in1=01010000 bcd_in2=10000001 cout=1 sum=00110001
* bcd_in1=01010000 bcd_in2=10000010 cout=1 sum=00110010
* bcd_in1=01010000 bcd_in2=10000011 cout=1 sum=00110011
* bcd_in1=01010000 bcd_in2=10000100 cout=1 sum=00110100
* bcd_in1=01010000 bcd_in2=10000101 cout=1 sum=00110101
* bcd_in1=01010000 bcd_in2=10000110 cout=1 sum=00110110
* bcd_in1=01010000 bcd_in2=10000111 cout=1 sum=00110111
* bcd_in1=01010000 bcd_in2=10001000 cout=1 sum=00111000
* bcd_in1=01010000 bcd_in2=10001001 cout=1 sum=00111001
* bcd_in1=01010000 bcd_in2=10010000 cout=1 sum=01000000
* bcd_in1=01010000 bcd_in2=10010001 cout=1 sum=01000001
* bcd_in1=01010000 bcd_in2=10010010 cout=1 sum=01000010
* bcd_in1=01010000 bcd_in2=10010011 cout=1 sum=01000011
* bcd_in1=01010000 bcd_in2=10010100 cout=1 sum=01000100
* bcd_in1=01010000 bcd_in2=10010101 cout=1 sum=01000101
* bcd_in1=01010000 bcd_in2=10010110 cout=1 sum=01000110
* bcd_in1=01010000 bcd_in2=10010111 cout=1 sum=01000111
* bcd_in1=01010000 bcd_in2=10011000 cout=1 sum=01001000
* bcd_in1=01010000 bcd_in2=10011001 cout=1 sum=01001001
* bcd_in1=01010001 bcd_in2=00000000 cout=0 sum=01010001
* bcd_in1=01010001 bcd_in2=00000001 cout=0 sum=01010010
* bcd_in1=01010001 bcd_in2=00000010 cout=0 sum=01010011
* bcd_in1=01010001 bcd_in2=00000011 cout=0 sum=01010100
* bcd_in1=01010001 bcd_in2=00000100 cout=0 sum=01010101
* bcd_in1=01010001 bcd_in2=00000101 cout=0 sum=01010110
* bcd_in1=01010001 bcd_in2=00000110 cout=0 sum=01010111
* bcd_in1=01010001 bcd_in2=00000111 cout=0 sum=01011000
* bcd_in1=01010001 bcd_in2=00001000 cout=0 sum=01011001
* bcd_in1=01010001 bcd_in2=00001001 cout=0 sum=01100000
* bcd_in1=01010001 bcd_in2=00010000 cout=0 sum=01100001
* bcd_in1=01010001 bcd_in2=00010001 cout=0 sum=01100010
* bcd_in1=01010001 bcd_in2=00010010 cout=0 sum=01100011
* bcd_in1=01010001 bcd_in2=00010011 cout=0 sum=01100100
* bcd_in1=01010001 bcd_in2=00010100 cout=0 sum=01100101
* bcd_in1=01010001 bcd_in2=00010101 cout=0 sum=01100110
* bcd_in1=01010001 bcd_in2=00010110 cout=0 sum=01100111
* bcd_in1=01010001 bcd_in2=00010111 cout=0 sum=01101000
* bcd_in1=01010001 bcd_in2=00011000 cout=0 sum=01101001
* bcd_in1=01010001 bcd_in2=00011001 cout=0 sum=01110000
* bcd_in1=01010001 bcd_in2=00100000 cout=0 sum=01110001
* bcd_in1=01010001 bcd_in2=00100001 cout=0 sum=01110010
* bcd_in1=01010001 bcd_in2=00100010 cout=0 sum=01110011
* bcd_in1=01010001 bcd_in2=00100011 cout=0 sum=01110100
* bcd_in1=01010001 bcd_in2=00100100 cout=0 sum=01110101
* bcd_in1=01010001 bcd_in2=00100101 cout=0 sum=01110110
* bcd_in1=01010001 bcd_in2=00100110 cout=0 sum=01110111
* bcd_in1=01010001 bcd_in2=00100111 cout=0 sum=01111000
* bcd_in1=01010001 bcd_in2=00101000 cout=0 sum=01111001
* bcd_in1=01010001 bcd_in2=00101001 cout=0 sum=10000000
* bcd_in1=01010001 bcd_in2=00110000 cout=0 sum=10000001
* bcd_in1=01010001 bcd_in2=00110001 cout=0 sum=10000010
* bcd_in1=01010001 bcd_in2=00110010 cout=0 sum=10000011
* bcd_in1=01010001 bcd_in2=00110011 cout=0 sum=10000100
* bcd_in1=01010001 bcd_in2=00110100 cout=0 sum=10000101
* bcd_in1=01010001 bcd_in2=00110101 cout=0 sum=10000110
* bcd_in1=01010001 bcd_in2=00110110 cout=0 sum=10000111
* bcd_in1=01010001 bcd_in2=00110111 cout=0 sum=10001000
* bcd_in1=01010001 bcd_in2=00111000 cout=0 sum=10001001
* bcd_in1=01010001 bcd_in2=00111001 cout=0 sum=10010000
* bcd_in1=01010001 bcd_in2=01000000 cout=0 sum=10010001
* bcd_in1=01010001 bcd_in2=01000001 cout=0 sum=10010010
* bcd_in1=01010001 bcd_in2=01000010 cout=0 sum=10010011
* bcd_in1=01010001 bcd_in2=01000011 cout=0 sum=10010100
* bcd_in1=01010001 bcd_in2=01000100 cout=0 sum=10010101
* bcd_in1=01010001 bcd_in2=01000101 cout=0 sum=10010110
* bcd_in1=01010001 bcd_in2=01000110 cout=0 sum=10010111
* bcd_in1=01010001 bcd_in2=01000111 cout=0 sum=10011000
* bcd_in1=01010001 bcd_in2=01001000 cout=0 sum=10011001
* bcd_in1=01010001 bcd_in2=01001001 cout=1 sum=00000000
* bcd_in1=01010001 bcd_in2=01010000 cout=1 sum=00000001
* bcd_in1=01010001 bcd_in2=01010001 cout=1 sum=00000010
* bcd_in1=01010001 bcd_in2=01010010 cout=1 sum=00000011
* bcd_in1=01010001 bcd_in2=01010011 cout=1 sum=00000100
* bcd_in1=01010001 bcd_in2=01010100 cout=1 sum=00000101
* bcd_in1=01010001 bcd_in2=01010101 cout=1 sum=00000110
* bcd_in1=01010001 bcd_in2=01010110 cout=1 sum=00000111
* bcd_in1=01010001 bcd_in2=01010111 cout=1 sum=00001000
* bcd_in1=01010001 bcd_in2=01011000 cout=1 sum=00001001
* bcd_in1=01010001 bcd_in2=01011001 cout=1 sum=00010000
* bcd_in1=01010001 bcd_in2=01100000 cout=1 sum=00010001
* bcd_in1=01010001 bcd_in2=01100001 cout=1 sum=00010010
* bcd_in1=01010001 bcd_in2=01100010 cout=1 sum=00010011
* bcd_in1=01010001 bcd_in2=01100011 cout=1 sum=00010100
* bcd_in1=01010001 bcd_in2=01100100 cout=1 sum=00010101
* bcd_in1=01010001 bcd_in2=01100101 cout=1 sum=00010110
* bcd_in1=01010001 bcd_in2=01100110 cout=1 sum=00010111
* bcd_in1=01010001 bcd_in2=01100111 cout=1 sum=00011000
* bcd_in1=01010001 bcd_in2=01101000 cout=1 sum=00011001
* bcd_in1=01010001 bcd_in2=01101001 cout=1 sum=00100000
* bcd_in1=01010001 bcd_in2=01110000 cout=1 sum=00100001
* bcd_in1=01010001 bcd_in2=01110001 cout=1 sum=00100010
* bcd_in1=01010001 bcd_in2=01110010 cout=1 sum=00100011
* bcd_in1=01010001 bcd_in2=01110011 cout=1 sum=00100100
* bcd_in1=01010001 bcd_in2=01110100 cout=1 sum=00100101
* bcd_in1=01010001 bcd_in2=01110101 cout=1 sum=00100110
* bcd_in1=01010001 bcd_in2=01110110 cout=1 sum=00100111
* bcd_in1=01010001 bcd_in2=01110111 cout=1 sum=00101000
* bcd_in1=01010001 bcd_in2=01111000 cout=1 sum=00101001
* bcd_in1=01010001 bcd_in2=01111001 cout=1 sum=00110000
* bcd_in1=01010001 bcd_in2=10000000 cout=1 sum=00110001
* bcd_in1=01010001 bcd_in2=10000001 cout=1 sum=00110010
* bcd_in1=01010001 bcd_in2=10000010 cout=1 sum=00110011
* bcd_in1=01010001 bcd_in2=10000011 cout=1 sum=00110100
* bcd_in1=01010001 bcd_in2=10000100 cout=1 sum=00110101
* bcd_in1=01010001 bcd_in2=10000101 cout=1 sum=00110110
* bcd_in1=01010001 bcd_in2=10000110 cout=1 sum=00110111
* bcd_in1=01010001 bcd_in2=10000111 cout=1 sum=00111000
* bcd_in1=01010001 bcd_in2=10001000 cout=1 sum=00111001
* bcd_in1=01010001 bcd_in2=10001001 cout=1 sum=01000000
* bcd_in1=01010001 bcd_in2=10010000 cout=1 sum=01000001
* bcd_in1=01010001 bcd_in2=10010001 cout=1 sum=01000010
* bcd_in1=01010001 bcd_in2=10010010 cout=1 sum=01000011
* bcd_in1=01010001 bcd_in2=10010011 cout=1 sum=01000100
* bcd_in1=01010001 bcd_in2=10010100 cout=1 sum=01000101
* bcd_in1=01010001 bcd_in2=10010101 cout=1 sum=01000110
* bcd_in1=01010001 bcd_in2=10010110 cout=1 sum=01000111
* bcd_in1=01010001 bcd_in2=10010111 cout=1 sum=01001000
* bcd_in1=01010001 bcd_in2=10011000 cout=1 sum=01001001
* bcd_in1=01010001 bcd_in2=10011001 cout=1 sum=01010000
* bcd_in1=01010010 bcd_in2=00000000 cout=0 sum=01010010
* bcd_in1=01010010 bcd_in2=00000001 cout=0 sum=01010011
* bcd_in1=01010010 bcd_in2=00000010 cout=0 sum=01010100
* bcd_in1=01010010 bcd_in2=00000011 cout=0 sum=01010101
* bcd_in1=01010010 bcd_in2=00000100 cout=0 sum=01010110
* bcd_in1=01010010 bcd_in2=00000101 cout=0 sum=01010111
* bcd_in1=01010010 bcd_in2=00000110 cout=0 sum=01011000
* bcd_in1=01010010 bcd_in2=00000111 cout=0 sum=01011001
* bcd_in1=01010010 bcd_in2=00001000 cout=0 sum=01100000
* bcd_in1=01010010 bcd_in2=00001001 cout=0 sum=01100001
* bcd_in1=01010010 bcd_in2=00010000 cout=0 sum=01100010
* bcd_in1=01010010 bcd_in2=00010001 cout=0 sum=01100011
* bcd_in1=01010010 bcd_in2=00010010 cout=0 sum=01100100
* bcd_in1=01010010 bcd_in2=00010011 cout=0 sum=01100101
* bcd_in1=01010010 bcd_in2=00010100 cout=0 sum=01100110
* bcd_in1=01010010 bcd_in2=00010101 cout=0 sum=01100111
* bcd_in1=01010010 bcd_in2=00010110 cout=0 sum=01101000
* bcd_in1=01010010 bcd_in2=00010111 cout=0 sum=01101001
* bcd_in1=01010010 bcd_in2=00011000 cout=0 sum=01110000
* bcd_in1=01010010 bcd_in2=00011001 cout=0 sum=01110001
* bcd_in1=01010010 bcd_in2=00100000 cout=0 sum=01110010
* bcd_in1=01010010 bcd_in2=00100001 cout=0 sum=01110011
* bcd_in1=01010010 bcd_in2=00100010 cout=0 sum=01110100
* bcd_in1=01010010 bcd_in2=00100011 cout=0 sum=01110101
* bcd_in1=01010010 bcd_in2=00100100 cout=0 sum=01110110
* bcd_in1=01010010 bcd_in2=00100101 cout=0 sum=01110111
* bcd_in1=01010010 bcd_in2=00100110 cout=0 sum=01111000
* bcd_in1=01010010 bcd_in2=00100111 cout=0 sum=01111001
* bcd_in1=01010010 bcd_in2=00101000 cout=0 sum=10000000
* bcd_in1=01010010 bcd_in2=00101001 cout=0 sum=10000001
* bcd_in1=01010010 bcd_in2=00110000 cout=0 sum=10000010
* bcd_in1=01010010 bcd_in2=00110001 cout=0 sum=10000011
* bcd_in1=01010010 bcd_in2=00110010 cout=0 sum=10000100
* bcd_in1=01010010 bcd_in2=00110011 cout=0 sum=10000101
* bcd_in1=01010010 bcd_in2=00110100 cout=0 sum=10000110
* bcd_in1=01010010 bcd_in2=00110101 cout=0 sum=10000111
* bcd_in1=01010010 bcd_in2=00110110 cout=0 sum=10001000
* bcd_in1=01010010 bcd_in2=00110111 cout=0 sum=10001001
* bcd_in1=01010010 bcd_in2=00111000 cout=0 sum=10010000
* bcd_in1=01010010 bcd_in2=00111001 cout=0 sum=10010001
* bcd_in1=01010010 bcd_in2=01000000 cout=0 sum=10010010
* bcd_in1=01010010 bcd_in2=01000001 cout=0 sum=10010011
* bcd_in1=01010010 bcd_in2=01000010 cout=0 sum=10010100
* bcd_in1=01010010 bcd_in2=01000011 cout=0 sum=10010101
* bcd_in1=01010010 bcd_in2=01000100 cout=0 sum=10010110
* bcd_in1=01010010 bcd_in2=01000101 cout=0 sum=10010111
* bcd_in1=01010010 bcd_in2=01000110 cout=0 sum=10011000
* bcd_in1=01010010 bcd_in2=01000111 cout=0 sum=10011001
* bcd_in1=01010010 bcd_in2=01001000 cout=1 sum=00000000
* bcd_in1=01010010 bcd_in2=01001001 cout=1 sum=00000001
* bcd_in1=01010010 bcd_in2=01010000 cout=1 sum=00000010
* bcd_in1=01010010 bcd_in2=01010001 cout=1 sum=00000011
* bcd_in1=01010010 bcd_in2=01010010 cout=1 sum=00000100
* bcd_in1=01010010 bcd_in2=01010011 cout=1 sum=00000101
* bcd_in1=01010010 bcd_in2=01010100 cout=1 sum=00000110
* bcd_in1=01010010 bcd_in2=01010101 cout=1 sum=00000111
* bcd_in1=01010010 bcd_in2=01010110 cout=1 sum=00001000
* bcd_in1=01010010 bcd_in2=01010111 cout=1 sum=00001001
* bcd_in1=01010010 bcd_in2=01011000 cout=1 sum=00010000
* bcd_in1=01010010 bcd_in2=01011001 cout=1 sum=00010001
* bcd_in1=01010010 bcd_in2=01100000 cout=1 sum=00010010
* bcd_in1=01010010 bcd_in2=01100001 cout=1 sum=00010011
* bcd_in1=01010010 bcd_in2=01100010 cout=1 sum=00010100
* bcd_in1=01010010 bcd_in2=01100011 cout=1 sum=00010101
* bcd_in1=01010010 bcd_in2=01100100 cout=1 sum=00010110
* bcd_in1=01010010 bcd_in2=01100101 cout=1 sum=00010111
* bcd_in1=01010010 bcd_in2=01100110 cout=1 sum=00011000
* bcd_in1=01010010 bcd_in2=01100111 cout=1 sum=00011001
* bcd_in1=01010010 bcd_in2=01101000 cout=1 sum=00100000
* bcd_in1=01010010 bcd_in2=01101001 cout=1 sum=00100001
* bcd_in1=01010010 bcd_in2=01110000 cout=1 sum=00100010
* bcd_in1=01010010 bcd_in2=01110001 cout=1 sum=00100011
* bcd_in1=01010010 bcd_in2=01110010 cout=1 sum=00100100
* bcd_in1=01010010 bcd_in2=01110011 cout=1 sum=00100101
* bcd_in1=01010010 bcd_in2=01110100 cout=1 sum=00100110
* bcd_in1=01010010 bcd_in2=01110101 cout=1 sum=00100111
* bcd_in1=01010010 bcd_in2=01110110 cout=1 sum=00101000
* bcd_in1=01010010 bcd_in2=01110111 cout=1 sum=00101001
* bcd_in1=01010010 bcd_in2=01111000 cout=1 sum=00110000
* bcd_in1=01010010 bcd_in2=01111001 cout=1 sum=00110001
* bcd_in1=01010010 bcd_in2=10000000 cout=1 sum=00110010
* bcd_in1=01010010 bcd_in2=10000001 cout=1 sum=00110011
* bcd_in1=01010010 bcd_in2=10000010 cout=1 sum=00110100
* bcd_in1=01010010 bcd_in2=10000011 cout=1 sum=00110101
* bcd_in1=01010010 bcd_in2=10000100 cout=1 sum=00110110
* bcd_in1=01010010 bcd_in2=10000101 cout=1 sum=00110111
* bcd_in1=01010010 bcd_in2=10000110 cout=1 sum=00111000
* bcd_in1=01010010 bcd_in2=10000111 cout=1 sum=00111001
* bcd_in1=01010010 bcd_in2=10001000 cout=1 sum=01000000
* bcd_in1=01010010 bcd_in2=10001001 cout=1 sum=01000001
* bcd_in1=01010010 bcd_in2=10010000 cout=1 sum=01000010
* bcd_in1=01010010 bcd_in2=10010001 cout=1 sum=01000011
* bcd_in1=01010010 bcd_in2=10010010 cout=1 sum=01000100
* bcd_in1=01010010 bcd_in2=10010011 cout=1 sum=01000101
* bcd_in1=01010010 bcd_in2=10010100 cout=1 sum=01000110
* bcd_in1=01010010 bcd_in2=10010101 cout=1 sum=01000111
* bcd_in1=01010010 bcd_in2=10010110 cout=1 sum=01001000
* bcd_in1=01010010 bcd_in2=10010111 cout=1 sum=01001001
* bcd_in1=01010010 bcd_in2=10011000 cout=1 sum=01010000
* bcd_in1=01010010 bcd_in2=10011001 cout=1 sum=01010001
* bcd_in1=01010011 bcd_in2=00000000 cout=0 sum=01010011
* bcd_in1=01010011 bcd_in2=00000001 cout=0 sum=01010100
* bcd_in1=01010011 bcd_in2=00000010 cout=0 sum=01010101
* bcd_in1=01010011 bcd_in2=00000011 cout=0 sum=01010110
* bcd_in1=01010011 bcd_in2=00000100 cout=0 sum=01010111
* bcd_in1=01010011 bcd_in2=00000101 cout=0 sum=01011000
* bcd_in1=01010011 bcd_in2=00000110 cout=0 sum=01011001
* bcd_in1=01010011 bcd_in2=00000111 cout=0 sum=01100000
* bcd_in1=01010011 bcd_in2=00001000 cout=0 sum=01100001
* bcd_in1=01010011 bcd_in2=00001001 cout=0 sum=01100010
* bcd_in1=01010011 bcd_in2=00010000 cout=0 sum=01100011
* bcd_in1=01010011 bcd_in2=00010001 cout=0 sum=01100100
* bcd_in1=01010011 bcd_in2=00010010 cout=0 sum=01100101
* bcd_in1=01010011 bcd_in2=00010011 cout=0 sum=01100110
* bcd_in1=01010011 bcd_in2=00010100 cout=0 sum=01100111
* bcd_in1=01010011 bcd_in2=00010101 cout=0 sum=01101000
* bcd_in1=01010011 bcd_in2=00010110 cout=0 sum=01101001
* bcd_in1=01010011 bcd_in2=00010111 cout=0 sum=01110000
* bcd_in1=01010011 bcd_in2=00011000 cout=0 sum=01110001
* bcd_in1=01010011 bcd_in2=00011001 cout=0 sum=01110010
* bcd_in1=01010011 bcd_in2=00100000 cout=0 sum=01110011
* bcd_in1=01010011 bcd_in2=00100001 cout=0 sum=01110100
* bcd_in1=01010011 bcd_in2=00100010 cout=0 sum=01110101
* bcd_in1=01010011 bcd_in2=00100011 cout=0 sum=01110110
* bcd_in1=01010011 bcd_in2=00100100 cout=0 sum=01110111
* bcd_in1=01010011 bcd_in2=00100101 cout=0 sum=01111000
* bcd_in1=01010011 bcd_in2=00100110 cout=0 sum=01111001
* bcd_in1=01010011 bcd_in2=00100111 cout=0 sum=10000000
* bcd_in1=01010011 bcd_in2=00101000 cout=0 sum=10000001
* bcd_in1=01010011 bcd_in2=00101001 cout=0 sum=10000010
* bcd_in1=01010011 bcd_in2=00110000 cout=0 sum=10000011
* bcd_in1=01010011 bcd_in2=00110001 cout=0 sum=10000100
* bcd_in1=01010011 bcd_in2=00110010 cout=0 sum=10000101
* bcd_in1=01010011 bcd_in2=00110011 cout=0 sum=10000110
* bcd_in1=01010011 bcd_in2=00110100 cout=0 sum=10000111
* bcd_in1=01010011 bcd_in2=00110101 cout=0 sum=10001000
* bcd_in1=01010011 bcd_in2=00110110 cout=0 sum=10001001
* bcd_in1=01010011 bcd_in2=00110111 cout=0 sum=10010000
* bcd_in1=01010011 bcd_in2=00111000 cout=0 sum=10010001
* bcd_in1=01010011 bcd_in2=00111001 cout=0 sum=10010010
* bcd_in1=01010011 bcd_in2=01000000 cout=0 sum=10010011
* bcd_in1=01010011 bcd_in2=01000001 cout=0 sum=10010100
* bcd_in1=01010011 bcd_in2=01000010 cout=0 sum=10010101
* bcd_in1=01010011 bcd_in2=01000011 cout=0 sum=10010110
* bcd_in1=01010011 bcd_in2=01000100 cout=0 sum=10010111
* bcd_in1=01010011 bcd_in2=01000101 cout=0 sum=10011000
* bcd_in1=01010011 bcd_in2=01000110 cout=0 sum=10011001
* bcd_in1=01010011 bcd_in2=01000111 cout=1 sum=00000000
* bcd_in1=01010011 bcd_in2=01001000 cout=1 sum=00000001
* bcd_in1=01010011 bcd_in2=01001001 cout=1 sum=00000010
* bcd_in1=01010011 bcd_in2=01010000 cout=1 sum=00000011
* bcd_in1=01010011 bcd_in2=01010001 cout=1 sum=00000100
* bcd_in1=01010011 bcd_in2=01010010 cout=1 sum=00000101
* bcd_in1=01010011 bcd_in2=01010011 cout=1 sum=00000110
* bcd_in1=01010011 bcd_in2=01010100 cout=1 sum=00000111
* bcd_in1=01010011 bcd_in2=01010101 cout=1 sum=00001000
* bcd_in1=01010011 bcd_in2=01010110 cout=1 sum=00001001
* bcd_in1=01010011 bcd_in2=01010111 cout=1 sum=00010000
* bcd_in1=01010011 bcd_in2=01011000 cout=1 sum=00010001
* bcd_in1=01010011 bcd_in2=01011001 cout=1 sum=00010010
* bcd_in1=01010011 bcd_in2=01100000 cout=1 sum=00010011
* bcd_in1=01010011 bcd_in2=01100001 cout=1 sum=00010100
* bcd_in1=01010011 bcd_in2=01100010 cout=1 sum=00010101
* bcd_in1=01010011 bcd_in2=01100011 cout=1 sum=00010110
* bcd_in1=01010011 bcd_in2=01100100 cout=1 sum=00010111
* bcd_in1=01010011 bcd_in2=01100101 cout=1 sum=00011000
* bcd_in1=01010011 bcd_in2=01100110 cout=1 sum=00011001
* bcd_in1=01010011 bcd_in2=01100111 cout=1 sum=00100000
* bcd_in1=01010011 bcd_in2=01101000 cout=1 sum=00100001
* bcd_in1=01010011 bcd_in2=01101001 cout=1 sum=00100010
* bcd_in1=01010011 bcd_in2=01110000 cout=1 sum=00100011
* bcd_in1=01010011 bcd_in2=01110001 cout=1 sum=00100100
* bcd_in1=01010011 bcd_in2=01110010 cout=1 sum=00100101
* bcd_in1=01010011 bcd_in2=01110011 cout=1 sum=00100110
* bcd_in1=01010011 bcd_in2=01110100 cout=1 sum=00100111
* bcd_in1=01010011 bcd_in2=01110101 cout=1 sum=00101000
* bcd_in1=01010011 bcd_in2=01110110 cout=1 sum=00101001
* bcd_in1=01010011 bcd_in2=01110111 cout=1 sum=00110000
* bcd_in1=01010011 bcd_in2=01111000 cout=1 sum=00110001
* bcd_in1=01010011 bcd_in2=01111001 cout=1 sum=00110010
* bcd_in1=01010011 bcd_in2=10000000 cout=1 sum=00110011
* bcd_in1=01010011 bcd_in2=10000001 cout=1 sum=00110100
* bcd_in1=01010011 bcd_in2=10000010 cout=1 sum=00110101
* bcd_in1=01010011 bcd_in2=10000011 cout=1 sum=00110110
* bcd_in1=01010011 bcd_in2=10000100 cout=1 sum=00110111
* bcd_in1=01010011 bcd_in2=10000101 cout=1 sum=00111000
* bcd_in1=01010011 bcd_in2=10000110 cout=1 sum=00111001
* bcd_in1=01010011 bcd_in2=10000111 cout=1 sum=01000000
* bcd_in1=01010011 bcd_in2=10001000 cout=1 sum=01000001
* bcd_in1=01010011 bcd_in2=10001001 cout=1 sum=01000010
* bcd_in1=01010011 bcd_in2=10010000 cout=1 sum=01000011
* bcd_in1=01010011 bcd_in2=10010001 cout=1 sum=01000100
* bcd_in1=01010011 bcd_in2=10010010 cout=1 sum=01000101
* bcd_in1=01010011 bcd_in2=10010011 cout=1 sum=01000110
* bcd_in1=01010011 bcd_in2=10010100 cout=1 sum=01000111
* bcd_in1=01010011 bcd_in2=10010101 cout=1 sum=01001000
* bcd_in1=01010011 bcd_in2=10010110 cout=1 sum=01001001
* bcd_in1=01010011 bcd_in2=10010111 cout=1 sum=01010000
* bcd_in1=01010011 bcd_in2=10011000 cout=1 sum=01010001
* bcd_in1=01010011 bcd_in2=10011001 cout=1 sum=01010010
* bcd_in1=01010100 bcd_in2=00000000 cout=0 sum=01010100
* bcd_in1=01010100 bcd_in2=00000001 cout=0 sum=01010101
* bcd_in1=01010100 bcd_in2=00000010 cout=0 sum=01010110
* bcd_in1=01010100 bcd_in2=00000011 cout=0 sum=01010111
* bcd_in1=01010100 bcd_in2=00000100 cout=0 sum=01011000
* bcd_in1=01010100 bcd_in2=00000101 cout=0 sum=01011001
* bcd_in1=01010100 bcd_in2=00000110 cout=0 sum=01100000
* bcd_in1=01010100 bcd_in2=00000111 cout=0 sum=01100001
* bcd_in1=01010100 bcd_in2=00001000 cout=0 sum=01100010
* bcd_in1=01010100 bcd_in2=00001001 cout=0 sum=01100011
* bcd_in1=01010100 bcd_in2=00010000 cout=0 sum=01100100
* bcd_in1=01010100 bcd_in2=00010001 cout=0 sum=01100101
* bcd_in1=01010100 bcd_in2=00010010 cout=0 sum=01100110
* bcd_in1=01010100 bcd_in2=00010011 cout=0 sum=01100111
* bcd_in1=01010100 bcd_in2=00010100 cout=0 sum=01101000
* bcd_in1=01010100 bcd_in2=00010101 cout=0 sum=01101001
* bcd_in1=01010100 bcd_in2=00010110 cout=0 sum=01110000
* bcd_in1=01010100 bcd_in2=00010111 cout=0 sum=01110001
* bcd_in1=01010100 bcd_in2=00011000 cout=0 sum=01110010
* bcd_in1=01010100 bcd_in2=00011001 cout=0 sum=01110011
* bcd_in1=01010100 bcd_in2=00100000 cout=0 sum=01110100
* bcd_in1=01010100 bcd_in2=00100001 cout=0 sum=01110101
* bcd_in1=01010100 bcd_in2=00100010 cout=0 sum=01110110
* bcd_in1=01010100 bcd_in2=00100011 cout=0 sum=01110111
* bcd_in1=01010100 bcd_in2=00100100 cout=0 sum=01111000
* bcd_in1=01010100 bcd_in2=00100101 cout=0 sum=01111001
* bcd_in1=01010100 bcd_in2=00100110 cout=0 sum=10000000
* bcd_in1=01010100 bcd_in2=00100111 cout=0 sum=10000001
* bcd_in1=01010100 bcd_in2=00101000 cout=0 sum=10000010
* bcd_in1=01010100 bcd_in2=00101001 cout=0 sum=10000011
* bcd_in1=01010100 bcd_in2=00110000 cout=0 sum=10000100
* bcd_in1=01010100 bcd_in2=00110001 cout=0 sum=10000101
* bcd_in1=01010100 bcd_in2=00110010 cout=0 sum=10000110
* bcd_in1=01010100 bcd_in2=00110011 cout=0 sum=10000111
* bcd_in1=01010100 bcd_in2=00110100 cout=0 sum=10001000
* bcd_in1=01010100 bcd_in2=00110101 cout=0 sum=10001001
* bcd_in1=01010100 bcd_in2=00110110 cout=0 sum=10010000
* bcd_in1=01010100 bcd_in2=00110111 cout=0 sum=10010001
* bcd_in1=01010100 bcd_in2=00111000 cout=0 sum=10010010
* bcd_in1=01010100 bcd_in2=00111001 cout=0 sum=10010011
* bcd_in1=01010100 bcd_in2=01000000 cout=0 sum=10010100
* bcd_in1=01010100 bcd_in2=01000001 cout=0 sum=10010101
* bcd_in1=01010100 bcd_in2=01000010 cout=0 sum=10010110
* bcd_in1=01010100 bcd_in2=01000011 cout=0 sum=10010111
* bcd_in1=01010100 bcd_in2=01000100 cout=0 sum=10011000
* bcd_in1=01010100 bcd_in2=01000101 cout=0 sum=10011001
* bcd_in1=01010100 bcd_in2=01000110 cout=1 sum=00000000
* bcd_in1=01010100 bcd_in2=01000111 cout=1 sum=00000001
* bcd_in1=01010100 bcd_in2=01001000 cout=1 sum=00000010
* bcd_in1=01010100 bcd_in2=01001001 cout=1 sum=00000011
* bcd_in1=01010100 bcd_in2=01010000 cout=1 sum=00000100
* bcd_in1=01010100 bcd_in2=01010001 cout=1 sum=00000101
* bcd_in1=01010100 bcd_in2=01010010 cout=1 sum=00000110
* bcd_in1=01010100 bcd_in2=01010011 cout=1 sum=00000111
* bcd_in1=01010100 bcd_in2=01010100 cout=1 sum=00001000
* bcd_in1=01010100 bcd_in2=01010101 cout=1 sum=00001001
* bcd_in1=01010100 bcd_in2=01010110 cout=1 sum=00010000
* bcd_in1=01010100 bcd_in2=01010111 cout=1 sum=00010001
* bcd_in1=01010100 bcd_in2=01011000 cout=1 sum=00010010
* bcd_in1=01010100 bcd_in2=01011001 cout=1 sum=00010011
* bcd_in1=01010100 bcd_in2=01100000 cout=1 sum=00010100
* bcd_in1=01010100 bcd_in2=01100001 cout=1 sum=00010101
* bcd_in1=01010100 bcd_in2=01100010 cout=1 sum=00010110
* bcd_in1=01010100 bcd_in2=01100011 cout=1 sum=00010111
* bcd_in1=01010100 bcd_in2=01100100 cout=1 sum=00011000
* bcd_in1=01010100 bcd_in2=01100101 cout=1 sum=00011001
* bcd_in1=01010100 bcd_in2=01100110 cout=1 sum=00100000
* bcd_in1=01010100 bcd_in2=01100111 cout=1 sum=00100001
* bcd_in1=01010100 bcd_in2=01101000 cout=1 sum=00100010
* bcd_in1=01010100 bcd_in2=01101001 cout=1 sum=00100011
* bcd_in1=01010100 bcd_in2=01110000 cout=1 sum=00100100
* bcd_in1=01010100 bcd_in2=01110001 cout=1 sum=00100101
* bcd_in1=01010100 bcd_in2=01110010 cout=1 sum=00100110
* bcd_in1=01010100 bcd_in2=01110011 cout=1 sum=00100111
* bcd_in1=01010100 bcd_in2=01110100 cout=1 sum=00101000
* bcd_in1=01010100 bcd_in2=01110101 cout=1 sum=00101001
* bcd_in1=01010100 bcd_in2=01110110 cout=1 sum=00110000
* bcd_in1=01010100 bcd_in2=01110111 cout=1 sum=00110001
* bcd_in1=01010100 bcd_in2=01111000 cout=1 sum=00110010
* bcd_in1=01010100 bcd_in2=01111001 cout=1 sum=00110011
* bcd_in1=01010100 bcd_in2=10000000 cout=1 sum=00110100
* bcd_in1=01010100 bcd_in2=10000001 cout=1 sum=00110101
* bcd_in1=01010100 bcd_in2=10000010 cout=1 sum=00110110
* bcd_in1=01010100 bcd_in2=10000011 cout=1 sum=00110111
* bcd_in1=01010100 bcd_in2=10000100 cout=1 sum=00111000
* bcd_in1=01010100 bcd_in2=10000101 cout=1 sum=00111001
* bcd_in1=01010100 bcd_in2=10000110 cout=1 sum=01000000
* bcd_in1=01010100 bcd_in2=10000111 cout=1 sum=01000001
* bcd_in1=01010100 bcd_in2=10001000 cout=1 sum=01000010
* bcd_in1=01010100 bcd_in2=10001001 cout=1 sum=01000011
* bcd_in1=01010100 bcd_in2=10010000 cout=1 sum=01000100
* bcd_in1=01010100 bcd_in2=10010001 cout=1 sum=01000101
* bcd_in1=01010100 bcd_in2=10010010 cout=1 sum=01000110
* bcd_in1=01010100 bcd_in2=10010011 cout=1 sum=01000111
* bcd_in1=01010100 bcd_in2=10010100 cout=1 sum=01001000
* bcd_in1=01010100 bcd_in2=10010101 cout=1 sum=01001001
* bcd_in1=01010100 bcd_in2=10010110 cout=1 sum=01010000
* bcd_in1=01010100 bcd_in2=10010111 cout=1 sum=01010001
* bcd_in1=01010100 bcd_in2=10011000 cout=1 sum=01010010
* bcd_in1=01010100 bcd_in2=10011001 cout=1 sum=01010011
* bcd_in1=01010101 bcd_in2=00000000 cout=0 sum=01010101
* bcd_in1=01010101 bcd_in2=00000001 cout=0 sum=01010110
* bcd_in1=01010101 bcd_in2=00000010 cout=0 sum=01010111
* bcd_in1=01010101 bcd_in2=00000011 cout=0 sum=01011000
* bcd_in1=01010101 bcd_in2=00000100 cout=0 sum=01011001
* bcd_in1=01010101 bcd_in2=00000101 cout=0 sum=01100000
* bcd_in1=01010101 bcd_in2=00000110 cout=0 sum=01100001
* bcd_in1=01010101 bcd_in2=00000111 cout=0 sum=01100010
* bcd_in1=01010101 bcd_in2=00001000 cout=0 sum=01100011
* bcd_in1=01010101 bcd_in2=00001001 cout=0 sum=01100100
* bcd_in1=01010101 bcd_in2=00010000 cout=0 sum=01100101
* bcd_in1=01010101 bcd_in2=00010001 cout=0 sum=01100110
* bcd_in1=01010101 bcd_in2=00010010 cout=0 sum=01100111
* bcd_in1=01010101 bcd_in2=00010011 cout=0 sum=01101000
* bcd_in1=01010101 bcd_in2=00010100 cout=0 sum=01101001
* bcd_in1=01010101 bcd_in2=00010101 cout=0 sum=01110000
* bcd_in1=01010101 bcd_in2=00010110 cout=0 sum=01110001
* bcd_in1=01010101 bcd_in2=00010111 cout=0 sum=01110010
* bcd_in1=01010101 bcd_in2=00011000 cout=0 sum=01110011
* bcd_in1=01010101 bcd_in2=00011001 cout=0 sum=01110100
* bcd_in1=01010101 bcd_in2=00100000 cout=0 sum=01110101
* bcd_in1=01010101 bcd_in2=00100001 cout=0 sum=01110110
* bcd_in1=01010101 bcd_in2=00100010 cout=0 sum=01110111
* bcd_in1=01010101 bcd_in2=00100011 cout=0 sum=01111000
* bcd_in1=01010101 bcd_in2=00100100 cout=0 sum=01111001
* bcd_in1=01010101 bcd_in2=00100101 cout=0 sum=10000000
* bcd_in1=01010101 bcd_in2=00100110 cout=0 sum=10000001
* bcd_in1=01010101 bcd_in2=00100111 cout=0 sum=10000010
* bcd_in1=01010101 bcd_in2=00101000 cout=0 sum=10000011
* bcd_in1=01010101 bcd_in2=00101001 cout=0 sum=10000100
* bcd_in1=01010101 bcd_in2=00110000 cout=0 sum=10000101
* bcd_in1=01010101 bcd_in2=00110001 cout=0 sum=10000110
* bcd_in1=01010101 bcd_in2=00110010 cout=0 sum=10000111
* bcd_in1=01010101 bcd_in2=00110011 cout=0 sum=10001000
* bcd_in1=01010101 bcd_in2=00110100 cout=0 sum=10001001
* bcd_in1=01010101 bcd_in2=00110101 cout=0 sum=10010000
* bcd_in1=01010101 bcd_in2=00110110 cout=0 sum=10010001
* bcd_in1=01010101 bcd_in2=00110111 cout=0 sum=10010010
* bcd_in1=01010101 bcd_in2=00111000 cout=0 sum=10010011
* bcd_in1=01010101 bcd_in2=00111001 cout=0 sum=10010100
* bcd_in1=01010101 bcd_in2=01000000 cout=0 sum=10010101
* bcd_in1=01010101 bcd_in2=01000001 cout=0 sum=10010110
* bcd_in1=01010101 bcd_in2=01000010 cout=0 sum=10010111
* bcd_in1=01010101 bcd_in2=01000011 cout=0 sum=10011000
* bcd_in1=01010101 bcd_in2=01000100 cout=0 sum=10011001
* bcd_in1=01010101 bcd_in2=01000101 cout=1 sum=00000000
* bcd_in1=01010101 bcd_in2=01000110 cout=1 sum=00000001
* bcd_in1=01010101 bcd_in2=01000111 cout=1 sum=00000010
* bcd_in1=01010101 bcd_in2=01001000 cout=1 sum=00000011
* bcd_in1=01010101 bcd_in2=01001001 cout=1 sum=00000100
* bcd_in1=01010101 bcd_in2=01010000 cout=1 sum=00000101
* bcd_in1=01010101 bcd_in2=01010001 cout=1 sum=00000110
* bcd_in1=01010101 bcd_in2=01010010 cout=1 sum=00000111
* bcd_in1=01010101 bcd_in2=01010011 cout=1 sum=00001000
* bcd_in1=01010101 bcd_in2=01010100 cout=1 sum=00001001
* bcd_in1=01010101 bcd_in2=01010101 cout=1 sum=00010000
* bcd_in1=01010101 bcd_in2=01010110 cout=1 sum=00010001
* bcd_in1=01010101 bcd_in2=01010111 cout=1 sum=00010010
* bcd_in1=01010101 bcd_in2=01011000 cout=1 sum=00010011
* bcd_in1=01010101 bcd_in2=01011001 cout=1 sum=00010100
* bcd_in1=01010101 bcd_in2=01100000 cout=1 sum=00010101
* bcd_in1=01010101 bcd_in2=01100001 cout=1 sum=00010110
* bcd_in1=01010101 bcd_in2=01100010 cout=1 sum=00010111
* bcd_in1=01010101 bcd_in2=01100011 cout=1 sum=00011000
* bcd_in1=01010101 bcd_in2=01100100 cout=1 sum=00011001
* bcd_in1=01010101 bcd_in2=01100101 cout=1 sum=00100000
* bcd_in1=01010101 bcd_in2=01100110 cout=1 sum=00100001
* bcd_in1=01010101 bcd_in2=01100111 cout=1 sum=00100010
* bcd_in1=01010101 bcd_in2=01101000 cout=1 sum=00100011
* bcd_in1=01010101 bcd_in2=01101001 cout=1 sum=00100100
* bcd_in1=01010101 bcd_in2=01110000 cout=1 sum=00100101
* bcd_in1=01010101 bcd_in2=01110001 cout=1 sum=00100110
* bcd_in1=01010101 bcd_in2=01110010 cout=1 sum=00100111
* bcd_in1=01010101 bcd_in2=01110011 cout=1 sum=00101000
* bcd_in1=01010101 bcd_in2=01110100 cout=1 sum=00101001
* bcd_in1=01010101 bcd_in2=01110101 cout=1 sum=00110000
* bcd_in1=01010101 bcd_in2=01110110 cout=1 sum=00110001
* bcd_in1=01010101 bcd_in2=01110111 cout=1 sum=00110010
* bcd_in1=01010101 bcd_in2=01111000 cout=1 sum=00110011
* bcd_in1=01010101 bcd_in2=01111001 cout=1 sum=00110100
* bcd_in1=01010101 bcd_in2=10000000 cout=1 sum=00110101
* bcd_in1=01010101 bcd_in2=10000001 cout=1 sum=00110110
* bcd_in1=01010101 bcd_in2=10000010 cout=1 sum=00110111
* bcd_in1=01010101 bcd_in2=10000011 cout=1 sum=00111000
* bcd_in1=01010101 bcd_in2=10000100 cout=1 sum=00111001
* bcd_in1=01010101 bcd_in2=10000101 cout=1 sum=01000000
* bcd_in1=01010101 bcd_in2=10000110 cout=1 sum=01000001
* bcd_in1=01010101 bcd_in2=10000111 cout=1 sum=01000010
* bcd_in1=01010101 bcd_in2=10001000 cout=1 sum=01000011
* bcd_in1=01010101 bcd_in2=10001001 cout=1 sum=01000100
* bcd_in1=01010101 bcd_in2=10010000 cout=1 sum=01000101
* bcd_in1=01010101 bcd_in2=10010001 cout=1 sum=01000110
* bcd_in1=01010101 bcd_in2=10010010 cout=1 sum=01000111
* bcd_in1=01010101 bcd_in2=10010011 cout=1 sum=01001000
* bcd_in1=01010101 bcd_in2=10010100 cout=1 sum=01001001
* bcd_in1=01010101 bcd_in2=10010101 cout=1 sum=01010000
* bcd_in1=01010101 bcd_in2=10010110 cout=1 sum=01010001
* bcd_in1=01010101 bcd_in2=10010111 cout=1 sum=01010010
* bcd_in1=01010101 bcd_in2=10011000 cout=1 sum=01010011
* bcd_in1=01010101 bcd_in2=10011001 cout=1 sum=01010100
* bcd_in1=01010110 bcd_in2=00000000 cout=0 sum=01010110
* bcd_in1=01010110 bcd_in2=00000001 cout=0 sum=01010111
* bcd_in1=01010110 bcd_in2=00000010 cout=0 sum=01011000
* bcd_in1=01010110 bcd_in2=00000011 cout=0 sum=01011001
* bcd_in1=01010110 bcd_in2=00000100 cout=0 sum=01100000
* bcd_in1=01010110 bcd_in2=00000101 cout=0 sum=01100001
* bcd_in1=01010110 bcd_in2=00000110 cout=0 sum=01100010
* bcd_in1=01010110 bcd_in2=00000111 cout=0 sum=01100011
* bcd_in1=01010110 bcd_in2=00001000 cout=0 sum=01100100
* bcd_in1=01010110 bcd_in2=00001001 cout=0 sum=01100101
* bcd_in1=01010110 bcd_in2=00010000 cout=0 sum=01100110
* bcd_in1=01010110 bcd_in2=00010001 cout=0 sum=01100111
* bcd_in1=01010110 bcd_in2=00010010 cout=0 sum=01101000
* bcd_in1=01010110 bcd_in2=00010011 cout=0 sum=01101001
* bcd_in1=01010110 bcd_in2=00010100 cout=0 sum=01110000
* bcd_in1=01010110 bcd_in2=00010101 cout=0 sum=01110001
* bcd_in1=01010110 bcd_in2=00010110 cout=0 sum=01110010
* bcd_in1=01010110 bcd_in2=00010111 cout=0 sum=01110011
* bcd_in1=01010110 bcd_in2=00011000 cout=0 sum=01110100
* bcd_in1=01010110 bcd_in2=00011001 cout=0 sum=01110101
* bcd_in1=01010110 bcd_in2=00100000 cout=0 sum=01110110
* bcd_in1=01010110 bcd_in2=00100001 cout=0 sum=01110111
* bcd_in1=01010110 bcd_in2=00100010 cout=0 sum=01111000
* bcd_in1=01010110 bcd_in2=00100011 cout=0 sum=01111001
* bcd_in1=01010110 bcd_in2=00100100 cout=0 sum=10000000
* bcd_in1=01010110 bcd_in2=00100101 cout=0 sum=10000001
* bcd_in1=01010110 bcd_in2=00100110 cout=0 sum=10000010
* bcd_in1=01010110 bcd_in2=00100111 cout=0 sum=10000011
* bcd_in1=01010110 bcd_in2=00101000 cout=0 sum=10000100
* bcd_in1=01010110 bcd_in2=00101001 cout=0 sum=10000101
* bcd_in1=01010110 bcd_in2=00110000 cout=0 sum=10000110
* bcd_in1=01010110 bcd_in2=00110001 cout=0 sum=10000111
* bcd_in1=01010110 bcd_in2=00110010 cout=0 sum=10001000
* bcd_in1=01010110 bcd_in2=00110011 cout=0 sum=10001001
* bcd_in1=01010110 bcd_in2=00110100 cout=0 sum=10010000
* bcd_in1=01010110 bcd_in2=00110101 cout=0 sum=10010001
* bcd_in1=01010110 bcd_in2=00110110 cout=0 sum=10010010
* bcd_in1=01010110 bcd_in2=00110111 cout=0 sum=10010011
* bcd_in1=01010110 bcd_in2=00111000 cout=0 sum=10010100
* bcd_in1=01010110 bcd_in2=00111001 cout=0 sum=10010101
* bcd_in1=01010110 bcd_in2=01000000 cout=0 sum=10010110
* bcd_in1=01010110 bcd_in2=01000001 cout=0 sum=10010111
* bcd_in1=01010110 bcd_in2=01000010 cout=0 sum=10011000
* bcd_in1=01010110 bcd_in2=01000011 cout=0 sum=10011001
* bcd_in1=01010110 bcd_in2=01000100 cout=1 sum=00000000
* bcd_in1=01010110 bcd_in2=01000101 cout=1 sum=00000001
* bcd_in1=01010110 bcd_in2=01000110 cout=1 sum=00000010
* bcd_in1=01010110 bcd_in2=01000111 cout=1 sum=00000011
* bcd_in1=01010110 bcd_in2=01001000 cout=1 sum=00000100
* bcd_in1=01010110 bcd_in2=01001001 cout=1 sum=00000101
* bcd_in1=01010110 bcd_in2=01010000 cout=1 sum=00000110
* bcd_in1=01010110 bcd_in2=01010001 cout=1 sum=00000111
* bcd_in1=01010110 bcd_in2=01010010 cout=1 sum=00001000
* bcd_in1=01010110 bcd_in2=01010011 cout=1 sum=00001001
* bcd_in1=01010110 bcd_in2=01010100 cout=1 sum=00010000
* bcd_in1=01010110 bcd_in2=01010101 cout=1 sum=00010001
* bcd_in1=01010110 bcd_in2=01010110 cout=1 sum=00010010
* bcd_in1=01010110 bcd_in2=01010111 cout=1 sum=00010011
* bcd_in1=01010110 bcd_in2=01011000 cout=1 sum=00010100
* bcd_in1=01010110 bcd_in2=01011001 cout=1 sum=00010101
* bcd_in1=01010110 bcd_in2=01100000 cout=1 sum=00010110
* bcd_in1=01010110 bcd_in2=01100001 cout=1 sum=00010111
* bcd_in1=01010110 bcd_in2=01100010 cout=1 sum=00011000
* bcd_in1=01010110 bcd_in2=01100011 cout=1 sum=00011001
* bcd_in1=01010110 bcd_in2=01100100 cout=1 sum=00100000
* bcd_in1=01010110 bcd_in2=01100101 cout=1 sum=00100001
* bcd_in1=01010110 bcd_in2=01100110 cout=1 sum=00100010
* bcd_in1=01010110 bcd_in2=01100111 cout=1 sum=00100011
* bcd_in1=01010110 bcd_in2=01101000 cout=1 sum=00100100
* bcd_in1=01010110 bcd_in2=01101001 cout=1 sum=00100101
* bcd_in1=01010110 bcd_in2=01110000 cout=1 sum=00100110
* bcd_in1=01010110 bcd_in2=01110001 cout=1 sum=00100111
* bcd_in1=01010110 bcd_in2=01110010 cout=1 sum=00101000
* bcd_in1=01010110 bcd_in2=01110011 cout=1 sum=00101001
* bcd_in1=01010110 bcd_in2=01110100 cout=1 sum=00110000
* bcd_in1=01010110 bcd_in2=01110101 cout=1 sum=00110001
* bcd_in1=01010110 bcd_in2=01110110 cout=1 sum=00110010
* bcd_in1=01010110 bcd_in2=01110111 cout=1 sum=00110011
* bcd_in1=01010110 bcd_in2=01111000 cout=1 sum=00110100
* bcd_in1=01010110 bcd_in2=01111001 cout=1 sum=00110101
* bcd_in1=01010110 bcd_in2=10000000 cout=1 sum=00110110
* bcd_in1=01010110 bcd_in2=10000001 cout=1 sum=00110111
* bcd_in1=01010110 bcd_in2=10000010 cout=1 sum=00111000
* bcd_in1=01010110 bcd_in2=10000011 cout=1 sum=00111001
* bcd_in1=01010110 bcd_in2=10000100 cout=1 sum=01000000
* bcd_in1=01010110 bcd_in2=10000101 cout=1 sum=01000001
* bcd_in1=01010110 bcd_in2=10000110 cout=1 sum=01000010
* bcd_in1=01010110 bcd_in2=10000111 cout=1 sum=01000011
* bcd_in1=01010110 bcd_in2=10001000 cout=1 sum=01000100
* bcd_in1=01010110 bcd_in2=10001001 cout=1 sum=01000101
* bcd_in1=01010110 bcd_in2=10010000 cout=1 sum=01000110
* bcd_in1=01010110 bcd_in2=10010001 cout=1 sum=01000111
* bcd_in1=01010110 bcd_in2=10010010 cout=1 sum=01001000
* bcd_in1=01010110 bcd_in2=10010011 cout=1 sum=01001001
* bcd_in1=01010110 bcd_in2=10010100 cout=1 sum=01010000
* bcd_in1=01010110 bcd_in2=10010101 cout=1 sum=01010001
* bcd_in1=01010110 bcd_in2=10010110 cout=1 sum=01010010
* bcd_in1=01010110 bcd_in2=10010111 cout=1 sum=01010011
* bcd_in1=01010110 bcd_in2=10011000 cout=1 sum=01010100
* bcd_in1=01010110 bcd_in2=10011001 cout=1 sum=01010101
* bcd_in1=01010111 bcd_in2=00000000 cout=0 sum=01010111
* bcd_in1=01010111 bcd_in2=00000001 cout=0 sum=01011000
* bcd_in1=01010111 bcd_in2=00000010 cout=0 sum=01011001
* bcd_in1=01010111 bcd_in2=00000011 cout=0 sum=01100000
* bcd_in1=01010111 bcd_in2=00000100 cout=0 sum=01100001
* bcd_in1=01010111 bcd_in2=00000101 cout=0 sum=01100010
* bcd_in1=01010111 bcd_in2=00000110 cout=0 sum=01100011
* bcd_in1=01010111 bcd_in2=00000111 cout=0 sum=01100100
* bcd_in1=01010111 bcd_in2=00001000 cout=0 sum=01100101
* bcd_in1=01010111 bcd_in2=00001001 cout=0 sum=01100110
* bcd_in1=01010111 bcd_in2=00010000 cout=0 sum=01100111
* bcd_in1=01010111 bcd_in2=00010001 cout=0 sum=01101000
* bcd_in1=01010111 bcd_in2=00010010 cout=0 sum=01101001
* bcd_in1=01010111 bcd_in2=00010011 cout=0 sum=01110000
* bcd_in1=01010111 bcd_in2=00010100 cout=0 sum=01110001
* bcd_in1=01010111 bcd_in2=00010101 cout=0 sum=01110010
* bcd_in1=01010111 bcd_in2=00010110 cout=0 sum=01110011
* bcd_in1=01010111 bcd_in2=00010111 cout=0 sum=01110100
* bcd_in1=01010111 bcd_in2=00011000 cout=0 sum=01110101
* bcd_in1=01010111 bcd_in2=00011001 cout=0 sum=01110110
* bcd_in1=01010111 bcd_in2=00100000 cout=0 sum=01110111
* bcd_in1=01010111 bcd_in2=00100001 cout=0 sum=01111000
* bcd_in1=01010111 bcd_in2=00100010 cout=0 sum=01111001
* bcd_in1=01010111 bcd_in2=00100011 cout=0 sum=10000000
* bcd_in1=01010111 bcd_in2=00100100 cout=0 sum=10000001
* bcd_in1=01010111 bcd_in2=00100101 cout=0 sum=10000010
* bcd_in1=01010111 bcd_in2=00100110 cout=0 sum=10000011
* bcd_in1=01010111 bcd_in2=00100111 cout=0 sum=10000100
* bcd_in1=01010111 bcd_in2=00101000 cout=0 sum=10000101
* bcd_in1=01010111 bcd_in2=00101001 cout=0 sum=10000110
* bcd_in1=01010111 bcd_in2=00110000 cout=0 sum=10000111
* bcd_in1=01010111 bcd_in2=00110001 cout=0 sum=10001000
* bcd_in1=01010111 bcd_in2=00110010 cout=0 sum=10001001
* bcd_in1=01010111 bcd_in2=00110011 cout=0 sum=10010000
* bcd_in1=01010111 bcd_in2=00110100 cout=0 sum=10010001
* bcd_in1=01010111 bcd_in2=00110101 cout=0 sum=10010010
* bcd_in1=01010111 bcd_in2=00110110 cout=0 sum=10010011
* bcd_in1=01010111 bcd_in2=00110111 cout=0 sum=10010100
* bcd_in1=01010111 bcd_in2=00111000 cout=0 sum=10010101
* bcd_in1=01010111 bcd_in2=00111001 cout=0 sum=10010110
* bcd_in1=01010111 bcd_in2=01000000 cout=0 sum=10010111
* bcd_in1=01010111 bcd_in2=01000001 cout=0 sum=10011000
* bcd_in1=01010111 bcd_in2=01000010 cout=0 sum=10011001
* bcd_in1=01010111 bcd_in2=01000011 cout=1 sum=00000000
* bcd_in1=01010111 bcd_in2=01000100 cout=1 sum=00000001
* bcd_in1=01010111 bcd_in2=01000101 cout=1 sum=00000010
* bcd_in1=01010111 bcd_in2=01000110 cout=1 sum=00000011
* bcd_in1=01010111 bcd_in2=01000111 cout=1 sum=00000100
* bcd_in1=01010111 bcd_in2=01001000 cout=1 sum=00000101
* bcd_in1=01010111 bcd_in2=01001001 cout=1 sum=00000110
* bcd_in1=01010111 bcd_in2=01010000 cout=1 sum=00000111
* bcd_in1=01010111 bcd_in2=01010001 cout=1 sum=00001000
* bcd_in1=01010111 bcd_in2=01010010 cout=1 sum=00001001
* bcd_in1=01010111 bcd_in2=01010011 cout=1 sum=00010000
* bcd_in1=01010111 bcd_in2=01010100 cout=1 sum=00010001
* bcd_in1=01010111 bcd_in2=01010101 cout=1 sum=00010010
* bcd_in1=01010111 bcd_in2=01010110 cout=1 sum=00010011
* bcd_in1=01010111 bcd_in2=01010111 cout=1 sum=00010100
* bcd_in1=01010111 bcd_in2=01011000 cout=1 sum=00010101
* bcd_in1=01010111 bcd_in2=01011001 cout=1 sum=00010110
* bcd_in1=01010111 bcd_in2=01100000 cout=1 sum=00010111
* bcd_in1=01010111 bcd_in2=01100001 cout=1 sum=00011000
* bcd_in1=01010111 bcd_in2=01100010 cout=1 sum=00011001
* bcd_in1=01010111 bcd_in2=01100011 cout=1 sum=00100000
* bcd_in1=01010111 bcd_in2=01100100 cout=1 sum=00100001
* bcd_in1=01010111 bcd_in2=01100101 cout=1 sum=00100010
* bcd_in1=01010111 bcd_in2=01100110 cout=1 sum=00100011
* bcd_in1=01010111 bcd_in2=01100111 cout=1 sum=00100100
* bcd_in1=01010111 bcd_in2=01101000 cout=1 sum=00100101
* bcd_in1=01010111 bcd_in2=01101001 cout=1 sum=00100110
* bcd_in1=01010111 bcd_in2=01110000 cout=1 sum=00100111
* bcd_in1=01010111 bcd_in2=01110001 cout=1 sum=00101000
* bcd_in1=01010111 bcd_in2=01110010 cout=1 sum=00101001
* bcd_in1=01010111 bcd_in2=01110011 cout=1 sum=00110000
* bcd_in1=01010111 bcd_in2=01110100 cout=1 sum=00110001
* bcd_in1=01010111 bcd_in2=01110101 cout=1 sum=00110010
* bcd_in1=01010111 bcd_in2=01110110 cout=1 sum=00110011
* bcd_in1=01010111 bcd_in2=01110111 cout=1 sum=00110100
* bcd_in1=01010111 bcd_in2=01111000 cout=1 sum=00110101
* bcd_in1=01010111 bcd_in2=01111001 cout=1 sum=00110110
* bcd_in1=01010111 bcd_in2=10000000 cout=1 sum=00110111
* bcd_in1=01010111 bcd_in2=10000001 cout=1 sum=00111000
* bcd_in1=01010111 bcd_in2=10000010 cout=1 sum=00111001
* bcd_in1=01010111 bcd_in2=10000011 cout=1 sum=01000000
* bcd_in1=01010111 bcd_in2=10000100 cout=1 sum=01000001
* bcd_in1=01010111 bcd_in2=10000101 cout=1 sum=01000010
* bcd_in1=01010111 bcd_in2=10000110 cout=1 sum=01000011
* bcd_in1=01010111 bcd_in2=10000111 cout=1 sum=01000100
* bcd_in1=01010111 bcd_in2=10001000 cout=1 sum=01000101
* bcd_in1=01010111 bcd_in2=10001001 cout=1 sum=01000110
* bcd_in1=01010111 bcd_in2=10010000 cout=1 sum=01000111
* bcd_in1=01010111 bcd_in2=10010001 cout=1 sum=01001000
* bcd_in1=01010111 bcd_in2=10010010 cout=1 sum=01001001
* bcd_in1=01010111 bcd_in2=10010011 cout=1 sum=01010000
* bcd_in1=01010111 bcd_in2=10010100 cout=1 sum=01010001
* bcd_in1=01010111 bcd_in2=10010101 cout=1 sum=01010010
* bcd_in1=01010111 bcd_in2=10010110 cout=1 sum=01010011
* bcd_in1=01010111 bcd_in2=10010111 cout=1 sum=01010100
* bcd_in1=01010111 bcd_in2=10011000 cout=1 sum=01010101
* bcd_in1=01010111 bcd_in2=10011001 cout=1 sum=01010110
* bcd_in1=01011000 bcd_in2=00000000 cout=0 sum=01011000
* bcd_in1=01011000 bcd_in2=00000001 cout=0 sum=01011001
* bcd_in1=01011000 bcd_in2=00000010 cout=0 sum=01100000
* bcd_in1=01011000 bcd_in2=00000011 cout=0 sum=01100001
* bcd_in1=01011000 bcd_in2=00000100 cout=0 sum=01100010
* bcd_in1=01011000 bcd_in2=00000101 cout=0 sum=01100011
* bcd_in1=01011000 bcd_in2=00000110 cout=0 sum=01100100
* bcd_in1=01011000 bcd_in2=00000111 cout=0 sum=01100101
* bcd_in1=01011000 bcd_in2=00001000 cout=0 sum=01100110
* bcd_in1=01011000 bcd_in2=00001001 cout=0 sum=01100111
* bcd_in1=01011000 bcd_in2=00010000 cout=0 sum=01101000
* bcd_in1=01011000 bcd_in2=00010001 cout=0 sum=01101001
* bcd_in1=01011000 bcd_in2=00010010 cout=0 sum=01110000
* bcd_in1=01011000 bcd_in2=00010011 cout=0 sum=01110001
* bcd_in1=01011000 bcd_in2=00010100 cout=0 sum=01110010
* bcd_in1=01011000 bcd_in2=00010101 cout=0 sum=01110011
* bcd_in1=01011000 bcd_in2=00010110 cout=0 sum=01110100
* bcd_in1=01011000 bcd_in2=00010111 cout=0 sum=01110101
* bcd_in1=01011000 bcd_in2=00011000 cout=0 sum=01110110
* bcd_in1=01011000 bcd_in2=00011001 cout=0 sum=01110111
* bcd_in1=01011000 bcd_in2=00100000 cout=0 sum=01111000
* bcd_in1=01011000 bcd_in2=00100001 cout=0 sum=01111001
* bcd_in1=01011000 bcd_in2=00100010 cout=0 sum=10000000
* bcd_in1=01011000 bcd_in2=00100011 cout=0 sum=10000001
* bcd_in1=01011000 bcd_in2=00100100 cout=0 sum=10000010
* bcd_in1=01011000 bcd_in2=00100101 cout=0 sum=10000011
* bcd_in1=01011000 bcd_in2=00100110 cout=0 sum=10000100
* bcd_in1=01011000 bcd_in2=00100111 cout=0 sum=10000101
* bcd_in1=01011000 bcd_in2=00101000 cout=0 sum=10000110
* bcd_in1=01011000 bcd_in2=00101001 cout=0 sum=10000111
* bcd_in1=01011000 bcd_in2=00110000 cout=0 sum=10001000
* bcd_in1=01011000 bcd_in2=00110001 cout=0 sum=10001001
* bcd_in1=01011000 bcd_in2=00110010 cout=0 sum=10010000
* bcd_in1=01011000 bcd_in2=00110011 cout=0 sum=10010001
* bcd_in1=01011000 bcd_in2=00110100 cout=0 sum=10010010
* bcd_in1=01011000 bcd_in2=00110101 cout=0 sum=10010011
* bcd_in1=01011000 bcd_in2=00110110 cout=0 sum=10010100
* bcd_in1=01011000 bcd_in2=00110111 cout=0 sum=10010101
* bcd_in1=01011000 bcd_in2=00111000 cout=0 sum=10010110
* bcd_in1=01011000 bcd_in2=00111001 cout=0 sum=10010111
* bcd_in1=01011000 bcd_in2=01000000 cout=0 sum=10011000
* bcd_in1=01011000 bcd_in2=01000001 cout=0 sum=10011001
* bcd_in1=01011000 bcd_in2=01000010 cout=1 sum=00000000
* bcd_in1=01011000 bcd_in2=01000011 cout=1 sum=00000001
* bcd_in1=01011000 bcd_in2=01000100 cout=1 sum=00000010
* bcd_in1=01011000 bcd_in2=01000101 cout=1 sum=00000011
* bcd_in1=01011000 bcd_in2=01000110 cout=1 sum=00000100
* bcd_in1=01011000 bcd_in2=01000111 cout=1 sum=00000101
* bcd_in1=01011000 bcd_in2=01001000 cout=1 sum=00000110
* bcd_in1=01011000 bcd_in2=01001001 cout=1 sum=00000111
* bcd_in1=01011000 bcd_in2=01010000 cout=1 sum=00001000
* bcd_in1=01011000 bcd_in2=01010001 cout=1 sum=00001001
* bcd_in1=01011000 bcd_in2=01010010 cout=1 sum=00010000
* bcd_in1=01011000 bcd_in2=01010011 cout=1 sum=00010001
* bcd_in1=01011000 bcd_in2=01010100 cout=1 sum=00010010
* bcd_in1=01011000 bcd_in2=01010101 cout=1 sum=00010011
* bcd_in1=01011000 bcd_in2=01010110 cout=1 sum=00010100
* bcd_in1=01011000 bcd_in2=01010111 cout=1 sum=00010101
* bcd_in1=01011000 bcd_in2=01011000 cout=1 sum=00010110
* bcd_in1=01011000 bcd_in2=01011001 cout=1 sum=00010111
* bcd_in1=01011000 bcd_in2=01100000 cout=1 sum=00011000
* bcd_in1=01011000 bcd_in2=01100001 cout=1 sum=00011001
* bcd_in1=01011000 bcd_in2=01100010 cout=1 sum=00100000
* bcd_in1=01011000 bcd_in2=01100011 cout=1 sum=00100001
* bcd_in1=01011000 bcd_in2=01100100 cout=1 sum=00100010
* bcd_in1=01011000 bcd_in2=01100101 cout=1 sum=00100011
* bcd_in1=01011000 bcd_in2=01100110 cout=1 sum=00100100
* bcd_in1=01011000 bcd_in2=01100111 cout=1 sum=00100101
* bcd_in1=01011000 bcd_in2=01101000 cout=1 sum=00100110
* bcd_in1=01011000 bcd_in2=01101001 cout=1 sum=00100111
* bcd_in1=01011000 bcd_in2=01110000 cout=1 sum=00101000
* bcd_in1=01011000 bcd_in2=01110001 cout=1 sum=00101001
* bcd_in1=01011000 bcd_in2=01110010 cout=1 sum=00110000
* bcd_in1=01011000 bcd_in2=01110011 cout=1 sum=00110001
* bcd_in1=01011000 bcd_in2=01110100 cout=1 sum=00110010
* bcd_in1=01011000 bcd_in2=01110101 cout=1 sum=00110011
* bcd_in1=01011000 bcd_in2=01110110 cout=1 sum=00110100
* bcd_in1=01011000 bcd_in2=01110111 cout=1 sum=00110101
* bcd_in1=01011000 bcd_in2=01111000 cout=1 sum=00110110
* bcd_in1=01011000 bcd_in2=01111001 cout=1 sum=00110111
* bcd_in1=01011000 bcd_in2=10000000 cout=1 sum=00111000
* bcd_in1=01011000 bcd_in2=10000001 cout=1 sum=00111001
* bcd_in1=01011000 bcd_in2=10000010 cout=1 sum=01000000
* bcd_in1=01011000 bcd_in2=10000011 cout=1 sum=01000001
* bcd_in1=01011000 bcd_in2=10000100 cout=1 sum=01000010
* bcd_in1=01011000 bcd_in2=10000101 cout=1 sum=01000011
* bcd_in1=01011000 bcd_in2=10000110 cout=1 sum=01000100
* bcd_in1=01011000 bcd_in2=10000111 cout=1 sum=01000101
* bcd_in1=01011000 bcd_in2=10001000 cout=1 sum=01000110
* bcd_in1=01011000 bcd_in2=10001001 cout=1 sum=01000111
* bcd_in1=01011000 bcd_in2=10010000 cout=1 sum=01001000
* bcd_in1=01011000 bcd_in2=10010001 cout=1 sum=01001001
* bcd_in1=01011000 bcd_in2=10010010 cout=1 sum=01010000
* bcd_in1=01011000 bcd_in2=10010011 cout=1 sum=01010001
* bcd_in1=01011000 bcd_in2=10010100 cout=1 sum=01010010
* bcd_in1=01011000 bcd_in2=10010101 cout=1 sum=01010011
* bcd_in1=01011000 bcd_in2=10010110 cout=1 sum=01010100
* bcd_in1=01011000 bcd_in2=10010111 cout=1 sum=01010101
* bcd_in1=01011000 bcd_in2=10011000 cout=1 sum=01010110
* bcd_in1=01011000 bcd_in2=10011001 cout=1 sum=01010111
* bcd_in1=01011001 bcd_in2=00000000 cout=0 sum=01011001
* bcd_in1=01011001 bcd_in2=00000001 cout=0 sum=01100000
* bcd_in1=01011001 bcd_in2=00000010 cout=0 sum=01100001
* bcd_in1=01011001 bcd_in2=00000011 cout=0 sum=01100010
* bcd_in1=01011001 bcd_in2=00000100 cout=0 sum=01100011
* bcd_in1=01011001 bcd_in2=00000101 cout=0 sum=01100100
* bcd_in1=01011001 bcd_in2=00000110 cout=0 sum=01100101
* bcd_in1=01011001 bcd_in2=00000111 cout=0 sum=01100110
* bcd_in1=01011001 bcd_in2=00001000 cout=0 sum=01100111
* bcd_in1=01011001 bcd_in2=00001001 cout=0 sum=01101000
* bcd_in1=01011001 bcd_in2=00010000 cout=0 sum=01101001
* bcd_in1=01011001 bcd_in2=00010001 cout=0 sum=01110000
* bcd_in1=01011001 bcd_in2=00010010 cout=0 sum=01110001
* bcd_in1=01011001 bcd_in2=00010011 cout=0 sum=01110010
* bcd_in1=01011001 bcd_in2=00010100 cout=0 sum=01110011
* bcd_in1=01011001 bcd_in2=00010101 cout=0 sum=01110100
* bcd_in1=01011001 bcd_in2=00010110 cout=0 sum=01110101
* bcd_in1=01011001 bcd_in2=00010111 cout=0 sum=01110110
* bcd_in1=01011001 bcd_in2=00011000 cout=0 sum=01110111
* bcd_in1=01011001 bcd_in2=00011001 cout=0 sum=01111000
* bcd_in1=01011001 bcd_in2=00100000 cout=0 sum=01111001
* bcd_in1=01011001 bcd_in2=00100001 cout=0 sum=10000000
* bcd_in1=01011001 bcd_in2=00100010 cout=0 sum=10000001
* bcd_in1=01011001 bcd_in2=00100011 cout=0 sum=10000010
* bcd_in1=01011001 bcd_in2=00100100 cout=0 sum=10000011
* bcd_in1=01011001 bcd_in2=00100101 cout=0 sum=10000100
* bcd_in1=01011001 bcd_in2=00100110 cout=0 sum=10000101
* bcd_in1=01011001 bcd_in2=00100111 cout=0 sum=10000110
* bcd_in1=01011001 bcd_in2=00101000 cout=0 sum=10000111
* bcd_in1=01011001 bcd_in2=00101001 cout=0 sum=10001000
* bcd_in1=01011001 bcd_in2=00110000 cout=0 sum=10001001
* bcd_in1=01011001 bcd_in2=00110001 cout=0 sum=10010000
* bcd_in1=01011001 bcd_in2=00110010 cout=0 sum=10010001
* bcd_in1=01011001 bcd_in2=00110011 cout=0 sum=10010010
* bcd_in1=01011001 bcd_in2=00110100 cout=0 sum=10010011
* bcd_in1=01011001 bcd_in2=00110101 cout=0 sum=10010100
* bcd_in1=01011001 bcd_in2=00110110 cout=0 sum=10010101
* bcd_in1=01011001 bcd_in2=00110111 cout=0 sum=10010110
* bcd_in1=01011001 bcd_in2=00111000 cout=0 sum=10010111
* bcd_in1=01011001 bcd_in2=00111001 cout=0 sum=10011000
* bcd_in1=01011001 bcd_in2=01000000 cout=0 sum=10011001
* bcd_in1=01011001 bcd_in2=01000001 cout=1 sum=00000000
* bcd_in1=01011001 bcd_in2=01000010 cout=1 sum=00000001
* bcd_in1=01011001 bcd_in2=01000011 cout=1 sum=00000010
* bcd_in1=01011001 bcd_in2=01000100 cout=1 sum=00000011
* bcd_in1=01011001 bcd_in2=01000101 cout=1 sum=00000100
* bcd_in1=01011001 bcd_in2=01000110 cout=1 sum=00000101
* bcd_in1=01011001 bcd_in2=01000111 cout=1 sum=00000110
* bcd_in1=01011001 bcd_in2=01001000 cout=1 sum=00000111
* bcd_in1=01011001 bcd_in2=01001001 cout=1 sum=00001000
* bcd_in1=01011001 bcd_in2=01010000 cout=1 sum=00001001
* bcd_in1=01011001 bcd_in2=01010001 cout=1 sum=00010000
* bcd_in1=01011001 bcd_in2=01010010 cout=1 sum=00010001
* bcd_in1=01011001 bcd_in2=01010011 cout=1 sum=00010010
* bcd_in1=01011001 bcd_in2=01010100 cout=1 sum=00010011
* bcd_in1=01011001 bcd_in2=01010101 cout=1 sum=00010100
* bcd_in1=01011001 bcd_in2=01010110 cout=1 sum=00010101
* bcd_in1=01011001 bcd_in2=01010111 cout=1 sum=00010110
* bcd_in1=01011001 bcd_in2=01011000 cout=1 sum=00010111
* bcd_in1=01011001 bcd_in2=01011001 cout=1 sum=00011000
* bcd_in1=01011001 bcd_in2=01100000 cout=1 sum=00011001
* bcd_in1=01011001 bcd_in2=01100001 cout=1 sum=00100000
* bcd_in1=01011001 bcd_in2=01100010 cout=1 sum=00100001
* bcd_in1=01011001 bcd_in2=01100011 cout=1 sum=00100010
* bcd_in1=01011001 bcd_in2=01100100 cout=1 sum=00100011
* bcd_in1=01011001 bcd_in2=01100101 cout=1 sum=00100100
* bcd_in1=01011001 bcd_in2=01100110 cout=1 sum=00100101
* bcd_in1=01011001 bcd_in2=01100111 cout=1 sum=00100110
* bcd_in1=01011001 bcd_in2=01101000 cout=1 sum=00100111
* bcd_in1=01011001 bcd_in2=01101001 cout=1 sum=00101000
* bcd_in1=01011001 bcd_in2=01110000 cout=1 sum=00101001
* bcd_in1=01011001 bcd_in2=01110001 cout=1 sum=00110000
* bcd_in1=01011001 bcd_in2=01110010 cout=1 sum=00110001
* bcd_in1=01011001 bcd_in2=01110011 cout=1 sum=00110010
* bcd_in1=01011001 bcd_in2=01110100 cout=1 sum=00110011
* bcd_in1=01011001 bcd_in2=01110101 cout=1 sum=00110100
* bcd_in1=01011001 bcd_in2=01110110 cout=1 sum=00110101
* bcd_in1=01011001 bcd_in2=01110111 cout=1 sum=00110110
* bcd_in1=01011001 bcd_in2=01111000 cout=1 sum=00110111
* bcd_in1=01011001 bcd_in2=01111001 cout=1 sum=00111000
* bcd_in1=01011001 bcd_in2=10000000 cout=1 sum=00111001
* bcd_in1=01011001 bcd_in2=10000001 cout=1 sum=01000000
* bcd_in1=01011001 bcd_in2=10000010 cout=1 sum=01000001
* bcd_in1=01011001 bcd_in2=10000011 cout=1 sum=01000010
* bcd_in1=01011001 bcd_in2=10000100 cout=1 sum=01000011
* bcd_in1=01011001 bcd_in2=10000101 cout=1 sum=01000100
* bcd_in1=01011001 bcd_in2=10000110 cout=1 sum=01000101
* bcd_in1=01011001 bcd_in2=10000111 cout=1 sum=01000110
* bcd_in1=01011001 bcd_in2=10001000 cout=1 sum=01000111
* bcd_in1=01011001 bcd_in2=10001001 cout=1 sum=01001000
* bcd_in1=01011001 bcd_in2=10010000 cout=1 sum=01001001
* bcd_in1=01011001 bcd_in2=10010001 cout=1 sum=01010000
* bcd_in1=01011001 bcd_in2=10010010 cout=1 sum=01010001
* bcd_in1=01011001 bcd_in2=10010011 cout=1 sum=01010010
* bcd_in1=01011001 bcd_in2=10010100 cout=1 sum=01010011
* bcd_in1=01011001 bcd_in2=10010101 cout=1 sum=01010100
* bcd_in1=01011001 bcd_in2=10010110 cout=1 sum=01010101
* bcd_in1=01011001 bcd_in2=10010111 cout=1 sum=01010110
* bcd_in1=01011001 bcd_in2=10011000 cout=1 sum=01010111
* bcd_in1=01011001 bcd_in2=10011001 cout=1 sum=01011000
* bcd_in1=01100000 bcd_in2=00000000 cout=0 sum=01100000
* bcd_in1=01100000 bcd_in2=00000001 cout=0 sum=01100001
* bcd_in1=01100000 bcd_in2=00000010 cout=0 sum=01100010
* bcd_in1=01100000 bcd_in2=00000011 cout=0 sum=01100011
* bcd_in1=01100000 bcd_in2=00000100 cout=0 sum=01100100
* bcd_in1=01100000 bcd_in2=00000101 cout=0 sum=01100101
* bcd_in1=01100000 bcd_in2=00000110 cout=0 sum=01100110
* bcd_in1=01100000 bcd_in2=00000111 cout=0 sum=01100111
* bcd_in1=01100000 bcd_in2=00001000 cout=0 sum=01101000
* bcd_in1=01100000 bcd_in2=00001001 cout=0 sum=01101001
* bcd_in1=01100000 bcd_in2=00010000 cout=0 sum=01110000
* bcd_in1=01100000 bcd_in2=00010001 cout=0 sum=01110001
* bcd_in1=01100000 bcd_in2=00010010 cout=0 sum=01110010
* bcd_in1=01100000 bcd_in2=00010011 cout=0 sum=01110011
* bcd_in1=01100000 bcd_in2=00010100 cout=0 sum=01110100
* bcd_in1=01100000 bcd_in2=00010101 cout=0 sum=01110101
* bcd_in1=01100000 bcd_in2=00010110 cout=0 sum=01110110
* bcd_in1=01100000 bcd_in2=00010111 cout=0 sum=01110111
* bcd_in1=01100000 bcd_in2=00011000 cout=0 sum=01111000
* bcd_in1=01100000 bcd_in2=00011001 cout=0 sum=01111001
* bcd_in1=01100000 bcd_in2=00100000 cout=0 sum=10000000
* bcd_in1=01100000 bcd_in2=00100001 cout=0 sum=10000001
* bcd_in1=01100000 bcd_in2=00100010 cout=0 sum=10000010
* bcd_in1=01100000 bcd_in2=00100011 cout=0 sum=10000011
* bcd_in1=01100000 bcd_in2=00100100 cout=0 sum=10000100
* bcd_in1=01100000 bcd_in2=00100101 cout=0 sum=10000101
* bcd_in1=01100000 bcd_in2=00100110 cout=0 sum=10000110
* bcd_in1=01100000 bcd_in2=00100111 cout=0 sum=10000111
* bcd_in1=01100000 bcd_in2=00101000 cout=0 sum=10001000
* bcd_in1=01100000 bcd_in2=00101001 cout=0 sum=10001001
* bcd_in1=01100000 bcd_in2=00110000 cout=0 sum=10010000
* bcd_in1=01100000 bcd_in2=00110001 cout=0 sum=10010001
* bcd_in1=01100000 bcd_in2=00110010 cout=0 sum=10010010
* bcd_in1=01100000 bcd_in2=00110011 cout=0 sum=10010011
* bcd_in1=01100000 bcd_in2=00110100 cout=0 sum=10010100
* bcd_in1=01100000 bcd_in2=00110101 cout=0 sum=10010101
* bcd_in1=01100000 bcd_in2=00110110 cout=0 sum=10010110
* bcd_in1=01100000 bcd_in2=00110111 cout=0 sum=10010111
* bcd_in1=01100000 bcd_in2=00111000 cout=0 sum=10011000
* bcd_in1=01100000 bcd_in2=00111001 cout=0 sum=10011001
* bcd_in1=01100000 bcd_in2=01000000 cout=1 sum=00000000
* bcd_in1=01100000 bcd_in2=01000001 cout=1 sum=00000001
* bcd_in1=01100000 bcd_in2=01000010 cout=1 sum=00000010
* bcd_in1=01100000 bcd_in2=01000011 cout=1 sum=00000011
* bcd_in1=01100000 bcd_in2=01000100 cout=1 sum=00000100
* bcd_in1=01100000 bcd_in2=01000101 cout=1 sum=00000101
* bcd_in1=01100000 bcd_in2=01000110 cout=1 sum=00000110
* bcd_in1=01100000 bcd_in2=01000111 cout=1 sum=00000111
* bcd_in1=01100000 bcd_in2=01001000 cout=1 sum=00001000
* bcd_in1=01100000 bcd_in2=01001001 cout=1 sum=00001001
* bcd_in1=01100000 bcd_in2=01010000 cout=1 sum=00010000
* bcd_in1=01100000 bcd_in2=01010001 cout=1 sum=00010001
* bcd_in1=01100000 bcd_in2=01010010 cout=1 sum=00010010
* bcd_in1=01100000 bcd_in2=01010011 cout=1 sum=00010011
* bcd_in1=01100000 bcd_in2=01010100 cout=1 sum=00010100
* bcd_in1=01100000 bcd_in2=01010101 cout=1 sum=00010101
* bcd_in1=01100000 bcd_in2=01010110 cout=1 sum=00010110
* bcd_in1=01100000 bcd_in2=01010111 cout=1 sum=00010111
* bcd_in1=01100000 bcd_in2=01011000 cout=1 sum=00011000
* bcd_in1=01100000 bcd_in2=01011001 cout=1 sum=00011001
* bcd_in1=01100000 bcd_in2=01100000 cout=1 sum=00100000
* bcd_in1=01100000 bcd_in2=01100001 cout=1 sum=00100001
* bcd_in1=01100000 bcd_in2=01100010 cout=1 sum=00100010
* bcd_in1=01100000 bcd_in2=01100011 cout=1 sum=00100011
* bcd_in1=01100000 bcd_in2=01100100 cout=1 sum=00100100
* bcd_in1=01100000 bcd_in2=01100101 cout=1 sum=00100101
* bcd_in1=01100000 bcd_in2=01100110 cout=1 sum=00100110
* bcd_in1=01100000 bcd_in2=01100111 cout=1 sum=00100111
* bcd_in1=01100000 bcd_in2=01101000 cout=1 sum=00101000
* bcd_in1=01100000 bcd_in2=01101001 cout=1 sum=00101001
* bcd_in1=01100000 bcd_in2=01110000 cout=1 sum=00110000
* bcd_in1=01100000 bcd_in2=01110001 cout=1 sum=00110001
* bcd_in1=01100000 bcd_in2=01110010 cout=1 sum=00110010
* bcd_in1=01100000 bcd_in2=01110011 cout=1 sum=00110011
* bcd_in1=01100000 bcd_in2=01110100 cout=1 sum=00110100
* bcd_in1=01100000 bcd_in2=01110101 cout=1 sum=00110101
* bcd_in1=01100000 bcd_in2=01110110 cout=1 sum=00110110
* bcd_in1=01100000 bcd_in2=01110111 cout=1 sum=00110111
* bcd_in1=01100000 bcd_in2=01111000 cout=1 sum=00111000
* bcd_in1=01100000 bcd_in2=01111001 cout=1 sum=00111001
* bcd_in1=01100000 bcd_in2=10000000 cout=1 sum=01000000
* bcd_in1=01100000 bcd_in2=10000001 cout=1 sum=01000001
* bcd_in1=01100000 bcd_in2=10000010 cout=1 sum=01000010
* bcd_in1=01100000 bcd_in2=10000011 cout=1 sum=01000011
* bcd_in1=01100000 bcd_in2=10000100 cout=1 sum=01000100
* bcd_in1=01100000 bcd_in2=10000101 cout=1 sum=01000101
* bcd_in1=01100000 bcd_in2=10000110 cout=1 sum=01000110
* bcd_in1=01100000 bcd_in2=10000111 cout=1 sum=01000111
* bcd_in1=01100000 bcd_in2=10001000 cout=1 sum=01001000
* bcd_in1=01100000 bcd_in2=10001001 cout=1 sum=01001001
* bcd_in1=01100000 bcd_in2=10010000 cout=1 sum=01010000
* bcd_in1=01100000 bcd_in2=10010001 cout=1 sum=01010001
* bcd_in1=01100000 bcd_in2=10010010 cout=1 sum=01010010
* bcd_in1=01100000 bcd_in2=10010011 cout=1 sum=01010011
* bcd_in1=01100000 bcd_in2=10010100 cout=1 sum=01010100
* bcd_in1=01100000 bcd_in2=10010101 cout=1 sum=01010101
* bcd_in1=01100000 bcd_in2=10010110 cout=1 sum=01010110
* bcd_in1=01100000 bcd_in2=10010111 cout=1 sum=01010111
* bcd_in1=01100000 bcd_in2=10011000 cout=1 sum=01011000
* bcd_in1=01100000 bcd_in2=10011001 cout=1 sum=01011001
* bcd_in1=01100001 bcd_in2=00000000 cout=0 sum=01100001
* bcd_in1=01100001 bcd_in2=00000001 cout=0 sum=01100010
* bcd_in1=01100001 bcd_in2=00000010 cout=0 sum=01100011
* bcd_in1=01100001 bcd_in2=00000011 cout=0 sum=01100100
* bcd_in1=01100001 bcd_in2=00000100 cout=0 sum=01100101
* bcd_in1=01100001 bcd_in2=00000101 cout=0 sum=01100110
* bcd_in1=01100001 bcd_in2=00000110 cout=0 sum=01100111
* bcd_in1=01100001 bcd_in2=00000111 cout=0 sum=01101000
* bcd_in1=01100001 bcd_in2=00001000 cout=0 sum=01101001
* bcd_in1=01100001 bcd_in2=00001001 cout=0 sum=01110000
* bcd_in1=01100001 bcd_in2=00010000 cout=0 sum=01110001
* bcd_in1=01100001 bcd_in2=00010001 cout=0 sum=01110010
* bcd_in1=01100001 bcd_in2=00010010 cout=0 sum=01110011
* bcd_in1=01100001 bcd_in2=00010011 cout=0 sum=01110100
* bcd_in1=01100001 bcd_in2=00010100 cout=0 sum=01110101
* bcd_in1=01100001 bcd_in2=00010101 cout=0 sum=01110110
* bcd_in1=01100001 bcd_in2=00010110 cout=0 sum=01110111
* bcd_in1=01100001 bcd_in2=00010111 cout=0 sum=01111000
* bcd_in1=01100001 bcd_in2=00011000 cout=0 sum=01111001
* bcd_in1=01100001 bcd_in2=00011001 cout=0 sum=10000000
* bcd_in1=01100001 bcd_in2=00100000 cout=0 sum=10000001
* bcd_in1=01100001 bcd_in2=00100001 cout=0 sum=10000010
* bcd_in1=01100001 bcd_in2=00100010 cout=0 sum=10000011
* bcd_in1=01100001 bcd_in2=00100011 cout=0 sum=10000100
* bcd_in1=01100001 bcd_in2=00100100 cout=0 sum=10000101
* bcd_in1=01100001 bcd_in2=00100101 cout=0 sum=10000110
* bcd_in1=01100001 bcd_in2=00100110 cout=0 sum=10000111
* bcd_in1=01100001 bcd_in2=00100111 cout=0 sum=10001000
* bcd_in1=01100001 bcd_in2=00101000 cout=0 sum=10001001
* bcd_in1=01100001 bcd_in2=00101001 cout=0 sum=10010000
* bcd_in1=01100001 bcd_in2=00110000 cout=0 sum=10010001
* bcd_in1=01100001 bcd_in2=00110001 cout=0 sum=10010010
* bcd_in1=01100001 bcd_in2=00110010 cout=0 sum=10010011
* bcd_in1=01100001 bcd_in2=00110011 cout=0 sum=10010100
* bcd_in1=01100001 bcd_in2=00110100 cout=0 sum=10010101
* bcd_in1=01100001 bcd_in2=00110101 cout=0 sum=10010110
* bcd_in1=01100001 bcd_in2=00110110 cout=0 sum=10010111
* bcd_in1=01100001 bcd_in2=00110111 cout=0 sum=10011000
* bcd_in1=01100001 bcd_in2=00111000 cout=0 sum=10011001
* bcd_in1=01100001 bcd_in2=00111001 cout=1 sum=00000000
* bcd_in1=01100001 bcd_in2=01000000 cout=1 sum=00000001
* bcd_in1=01100001 bcd_in2=01000001 cout=1 sum=00000010
* bcd_in1=01100001 bcd_in2=01000010 cout=1 sum=00000011
* bcd_in1=01100001 bcd_in2=01000011 cout=1 sum=00000100
* bcd_in1=01100001 bcd_in2=01000100 cout=1 sum=00000101
* bcd_in1=01100001 bcd_in2=01000101 cout=1 sum=00000110
* bcd_in1=01100001 bcd_in2=01000110 cout=1 sum=00000111
* bcd_in1=01100001 bcd_in2=01000111 cout=1 sum=00001000
* bcd_in1=01100001 bcd_in2=01001000 cout=1 sum=00001001
* bcd_in1=01100001 bcd_in2=01001001 cout=1 sum=00010000
* bcd_in1=01100001 bcd_in2=01010000 cout=1 sum=00010001
* bcd_in1=01100001 bcd_in2=01010001 cout=1 sum=00010010
* bcd_in1=01100001 bcd_in2=01010010 cout=1 sum=00010011
* bcd_in1=01100001 bcd_in2=01010011 cout=1 sum=00010100
* bcd_in1=01100001 bcd_in2=01010100 cout=1 sum=00010101
* bcd_in1=01100001 bcd_in2=01010101 cout=1 sum=00010110
* bcd_in1=01100001 bcd_in2=01010110 cout=1 sum=00010111
* bcd_in1=01100001 bcd_in2=01010111 cout=1 sum=00011000
* bcd_in1=01100001 bcd_in2=01011000 cout=1 sum=00011001
* bcd_in1=01100001 bcd_in2=01011001 cout=1 sum=00100000
* bcd_in1=01100001 bcd_in2=01100000 cout=1 sum=00100001
* bcd_in1=01100001 bcd_in2=01100001 cout=1 sum=00100010
* bcd_in1=01100001 bcd_in2=01100010 cout=1 sum=00100011
* bcd_in1=01100001 bcd_in2=01100011 cout=1 sum=00100100
* bcd_in1=01100001 bcd_in2=01100100 cout=1 sum=00100101
* bcd_in1=01100001 bcd_in2=01100101 cout=1 sum=00100110
* bcd_in1=01100001 bcd_in2=01100110 cout=1 sum=00100111
* bcd_in1=01100001 bcd_in2=01100111 cout=1 sum=00101000
* bcd_in1=01100001 bcd_in2=01101000 cout=1 sum=00101001
* bcd_in1=01100001 bcd_in2=01101001 cout=1 sum=00110000
* bcd_in1=01100001 bcd_in2=01110000 cout=1 sum=00110001
* bcd_in1=01100001 bcd_in2=01110001 cout=1 sum=00110010
* bcd_in1=01100001 bcd_in2=01110010 cout=1 sum=00110011
* bcd_in1=01100001 bcd_in2=01110011 cout=1 sum=00110100
* bcd_in1=01100001 bcd_in2=01110100 cout=1 sum=00110101
* bcd_in1=01100001 bcd_in2=01110101 cout=1 sum=00110110
* bcd_in1=01100001 bcd_in2=01110110 cout=1 sum=00110111
* bcd_in1=01100001 bcd_in2=01110111 cout=1 sum=00111000
* bcd_in1=01100001 bcd_in2=01111000 cout=1 sum=00111001
* bcd_in1=01100001 bcd_in2=01111001 cout=1 sum=01000000
* bcd_in1=01100001 bcd_in2=10000000 cout=1 sum=01000001
* bcd_in1=01100001 bcd_in2=10000001 cout=1 sum=01000010
* bcd_in1=01100001 bcd_in2=10000010 cout=1 sum=01000011
* bcd_in1=01100001 bcd_in2=10000011 cout=1 sum=01000100
* bcd_in1=01100001 bcd_in2=10000100 cout=1 sum=01000101
* bcd_in1=01100001 bcd_in2=10000101 cout=1 sum=01000110
* bcd_in1=01100001 bcd_in2=10000110 cout=1 sum=01000111
* bcd_in1=01100001 bcd_in2=10000111 cout=1 sum=01001000
* bcd_in1=01100001 bcd_in2=10001000 cout=1 sum=01001001
* bcd_in1=01100001 bcd_in2=10001001 cout=1 sum=01010000
* bcd_in1=01100001 bcd_in2=10010000 cout=1 sum=01010001
* bcd_in1=01100001 bcd_in2=10010001 cout=1 sum=01010010
* bcd_in1=01100001 bcd_in2=10010010 cout=1 sum=01010011
* bcd_in1=01100001 bcd_in2=10010011 cout=1 sum=01010100
* bcd_in1=01100001 bcd_in2=10010100 cout=1 sum=01010101
* bcd_in1=01100001 bcd_in2=10010101 cout=1 sum=01010110
* bcd_in1=01100001 bcd_in2=10010110 cout=1 sum=01010111
* bcd_in1=01100001 bcd_in2=10010111 cout=1 sum=01011000
* bcd_in1=01100001 bcd_in2=10011000 cout=1 sum=01011001
* bcd_in1=01100001 bcd_in2=10011001 cout=1 sum=01100000
* bcd_in1=01100010 bcd_in2=00000000 cout=0 sum=01100010
* bcd_in1=01100010 bcd_in2=00000001 cout=0 sum=01100011
* bcd_in1=01100010 bcd_in2=00000010 cout=0 sum=01100100
* bcd_in1=01100010 bcd_in2=00000011 cout=0 sum=01100101
* bcd_in1=01100010 bcd_in2=00000100 cout=0 sum=01100110
* bcd_in1=01100010 bcd_in2=00000101 cout=0 sum=01100111
* bcd_in1=01100010 bcd_in2=00000110 cout=0 sum=01101000
* bcd_in1=01100010 bcd_in2=00000111 cout=0 sum=01101001
* bcd_in1=01100010 bcd_in2=00001000 cout=0 sum=01110000
* bcd_in1=01100010 bcd_in2=00001001 cout=0 sum=01110001
* bcd_in1=01100010 bcd_in2=00010000 cout=0 sum=01110010
* bcd_in1=01100010 bcd_in2=00010001 cout=0 sum=01110011
* bcd_in1=01100010 bcd_in2=00010010 cout=0 sum=01110100
* bcd_in1=01100010 bcd_in2=00010011 cout=0 sum=01110101
* bcd_in1=01100010 bcd_in2=00010100 cout=0 sum=01110110
* bcd_in1=01100010 bcd_in2=00010101 cout=0 sum=01110111
* bcd_in1=01100010 bcd_in2=00010110 cout=0 sum=01111000
* bcd_in1=01100010 bcd_in2=00010111 cout=0 sum=01111001
* bcd_in1=01100010 bcd_in2=00011000 cout=0 sum=10000000
* bcd_in1=01100010 bcd_in2=00011001 cout=0 sum=10000001
* bcd_in1=01100010 bcd_in2=00100000 cout=0 sum=10000010
* bcd_in1=01100010 bcd_in2=00100001 cout=0 sum=10000011
* bcd_in1=01100010 bcd_in2=00100010 cout=0 sum=10000100
* bcd_in1=01100010 bcd_in2=00100011 cout=0 sum=10000101
* bcd_in1=01100010 bcd_in2=00100100 cout=0 sum=10000110
* bcd_in1=01100010 bcd_in2=00100101 cout=0 sum=10000111
* bcd_in1=01100010 bcd_in2=00100110 cout=0 sum=10001000
* bcd_in1=01100010 bcd_in2=00100111 cout=0 sum=10001001
* bcd_in1=01100010 bcd_in2=00101000 cout=0 sum=10010000
* bcd_in1=01100010 bcd_in2=00101001 cout=0 sum=10010001
* bcd_in1=01100010 bcd_in2=00110000 cout=0 sum=10010010
* bcd_in1=01100010 bcd_in2=00110001 cout=0 sum=10010011
* bcd_in1=01100010 bcd_in2=00110010 cout=0 sum=10010100
* bcd_in1=01100010 bcd_in2=00110011 cout=0 sum=10010101
* bcd_in1=01100010 bcd_in2=00110100 cout=0 sum=10010110
* bcd_in1=01100010 bcd_in2=00110101 cout=0 sum=10010111
* bcd_in1=01100010 bcd_in2=00110110 cout=0 sum=10011000
* bcd_in1=01100010 bcd_in2=00110111 cout=0 sum=10011001
* bcd_in1=01100010 bcd_in2=00111000 cout=1 sum=00000000
* bcd_in1=01100010 bcd_in2=00111001 cout=1 sum=00000001
* bcd_in1=01100010 bcd_in2=01000000 cout=1 sum=00000010
* bcd_in1=01100010 bcd_in2=01000001 cout=1 sum=00000011
* bcd_in1=01100010 bcd_in2=01000010 cout=1 sum=00000100
* bcd_in1=01100010 bcd_in2=01000011 cout=1 sum=00000101
* bcd_in1=01100010 bcd_in2=01000100 cout=1 sum=00000110
* bcd_in1=01100010 bcd_in2=01000101 cout=1 sum=00000111
* bcd_in1=01100010 bcd_in2=01000110 cout=1 sum=00001000
* bcd_in1=01100010 bcd_in2=01000111 cout=1 sum=00001001
* bcd_in1=01100010 bcd_in2=01001000 cout=1 sum=00010000
* bcd_in1=01100010 bcd_in2=01001001 cout=1 sum=00010001
* bcd_in1=01100010 bcd_in2=01010000 cout=1 sum=00010010
* bcd_in1=01100010 bcd_in2=01010001 cout=1 sum=00010011
* bcd_in1=01100010 bcd_in2=01010010 cout=1 sum=00010100
* bcd_in1=01100010 bcd_in2=01010011 cout=1 sum=00010101
* bcd_in1=01100010 bcd_in2=01010100 cout=1 sum=00010110
* bcd_in1=01100010 bcd_in2=01010101 cout=1 sum=00010111
* bcd_in1=01100010 bcd_in2=01010110 cout=1 sum=00011000
* bcd_in1=01100010 bcd_in2=01010111 cout=1 sum=00011001
* bcd_in1=01100010 bcd_in2=01011000 cout=1 sum=00100000
* bcd_in1=01100010 bcd_in2=01011001 cout=1 sum=00100001
* bcd_in1=01100010 bcd_in2=01100000 cout=1 sum=00100010
* bcd_in1=01100010 bcd_in2=01100001 cout=1 sum=00100011
* bcd_in1=01100010 bcd_in2=01100010 cout=1 sum=00100100
* bcd_in1=01100010 bcd_in2=01100011 cout=1 sum=00100101
* bcd_in1=01100010 bcd_in2=01100100 cout=1 sum=00100110
* bcd_in1=01100010 bcd_in2=01100101 cout=1 sum=00100111
* bcd_in1=01100010 bcd_in2=01100110 cout=1 sum=00101000
* bcd_in1=01100010 bcd_in2=01100111 cout=1 sum=00101001
* bcd_in1=01100010 bcd_in2=01101000 cout=1 sum=00110000
* bcd_in1=01100010 bcd_in2=01101001 cout=1 sum=00110001
* bcd_in1=01100010 bcd_in2=01110000 cout=1 sum=00110010
* bcd_in1=01100010 bcd_in2=01110001 cout=1 sum=00110011
* bcd_in1=01100010 bcd_in2=01110010 cout=1 sum=00110100
* bcd_in1=01100010 bcd_in2=01110011 cout=1 sum=00110101
* bcd_in1=01100010 bcd_in2=01110100 cout=1 sum=00110110
* bcd_in1=01100010 bcd_in2=01110101 cout=1 sum=00110111
* bcd_in1=01100010 bcd_in2=01110110 cout=1 sum=00111000
* bcd_in1=01100010 bcd_in2=01110111 cout=1 sum=00111001
* bcd_in1=01100010 bcd_in2=01111000 cout=1 sum=01000000
* bcd_in1=01100010 bcd_in2=01111001 cout=1 sum=01000001
* bcd_in1=01100010 bcd_in2=10000000 cout=1 sum=01000010
* bcd_in1=01100010 bcd_in2=10000001 cout=1 sum=01000011
* bcd_in1=01100010 bcd_in2=10000010 cout=1 sum=01000100
* bcd_in1=01100010 bcd_in2=10000011 cout=1 sum=01000101
* bcd_in1=01100010 bcd_in2=10000100 cout=1 sum=01000110
* bcd_in1=01100010 bcd_in2=10000101 cout=1 sum=01000111
* bcd_in1=01100010 bcd_in2=10000110 cout=1 sum=01001000
* bcd_in1=01100010 bcd_in2=10000111 cout=1 sum=01001001
* bcd_in1=01100010 bcd_in2=10001000 cout=1 sum=01010000
* bcd_in1=01100010 bcd_in2=10001001 cout=1 sum=01010001
* bcd_in1=01100010 bcd_in2=10010000 cout=1 sum=01010010
* bcd_in1=01100010 bcd_in2=10010001 cout=1 sum=01010011
* bcd_in1=01100010 bcd_in2=10010010 cout=1 sum=01010100
* bcd_in1=01100010 bcd_in2=10010011 cout=1 sum=01010101
* bcd_in1=01100010 bcd_in2=10010100 cout=1 sum=01010110
* bcd_in1=01100010 bcd_in2=10010101 cout=1 sum=01010111
* bcd_in1=01100010 bcd_in2=10010110 cout=1 sum=01011000
* bcd_in1=01100010 bcd_in2=10010111 cout=1 sum=01011001
* bcd_in1=01100010 bcd_in2=10011000 cout=1 sum=01100000
* bcd_in1=01100010 bcd_in2=10011001 cout=1 sum=01100001
* bcd_in1=01100011 bcd_in2=00000000 cout=0 sum=01100011
* bcd_in1=01100011 bcd_in2=00000001 cout=0 sum=01100100
* bcd_in1=01100011 bcd_in2=00000010 cout=0 sum=01100101
* bcd_in1=01100011 bcd_in2=00000011 cout=0 sum=01100110
* bcd_in1=01100011 bcd_in2=00000100 cout=0 sum=01100111
* bcd_in1=01100011 bcd_in2=00000101 cout=0 sum=01101000
* bcd_in1=01100011 bcd_in2=00000110 cout=0 sum=01101001
* bcd_in1=01100011 bcd_in2=00000111 cout=0 sum=01110000
* bcd_in1=01100011 bcd_in2=00001000 cout=0 sum=01110001
* bcd_in1=01100011 bcd_in2=00001001 cout=0 sum=01110010
* bcd_in1=01100011 bcd_in2=00010000 cout=0 sum=01110011
* bcd_in1=01100011 bcd_in2=00010001 cout=0 sum=01110100
* bcd_in1=01100011 bcd_in2=00010010 cout=0 sum=01110101
* bcd_in1=01100011 bcd_in2=00010011 cout=0 sum=01110110
* bcd_in1=01100011 bcd_in2=00010100 cout=0 sum=01110111
* bcd_in1=01100011 bcd_in2=00010101 cout=0 sum=01111000
* bcd_in1=01100011 bcd_in2=00010110 cout=0 sum=01111001
* bcd_in1=01100011 bcd_in2=00010111 cout=0 sum=10000000
* bcd_in1=01100011 bcd_in2=00011000 cout=0 sum=10000001
* bcd_in1=01100011 bcd_in2=00011001 cout=0 sum=10000010
* bcd_in1=01100011 bcd_in2=00100000 cout=0 sum=10000011
* bcd_in1=01100011 bcd_in2=00100001 cout=0 sum=10000100
* bcd_in1=01100011 bcd_in2=00100010 cout=0 sum=10000101
* bcd_in1=01100011 bcd_in2=00100011 cout=0 sum=10000110
* bcd_in1=01100011 bcd_in2=00100100 cout=0 sum=10000111
* bcd_in1=01100011 bcd_in2=00100101 cout=0 sum=10001000
* bcd_in1=01100011 bcd_in2=00100110 cout=0 sum=10001001
* bcd_in1=01100011 bcd_in2=00100111 cout=0 sum=10010000
* bcd_in1=01100011 bcd_in2=00101000 cout=0 sum=10010001
* bcd_in1=01100011 bcd_in2=00101001 cout=0 sum=10010010
* bcd_in1=01100011 bcd_in2=00110000 cout=0 sum=10010011
* bcd_in1=01100011 bcd_in2=00110001 cout=0 sum=10010100
* bcd_in1=01100011 bcd_in2=00110010 cout=0 sum=10010101
* bcd_in1=01100011 bcd_in2=00110011 cout=0 sum=10010110
* bcd_in1=01100011 bcd_in2=00110100 cout=0 sum=10010111
* bcd_in1=01100011 bcd_in2=00110101 cout=0 sum=10011000
* bcd_in1=01100011 bcd_in2=00110110 cout=0 sum=10011001
* bcd_in1=01100011 bcd_in2=00110111 cout=1 sum=00000000
* bcd_in1=01100011 bcd_in2=00111000 cout=1 sum=00000001
* bcd_in1=01100011 bcd_in2=00111001 cout=1 sum=00000010
* bcd_in1=01100011 bcd_in2=01000000 cout=1 sum=00000011
* bcd_in1=01100011 bcd_in2=01000001 cout=1 sum=00000100
* bcd_in1=01100011 bcd_in2=01000010 cout=1 sum=00000101
* bcd_in1=01100011 bcd_in2=01000011 cout=1 sum=00000110
* bcd_in1=01100011 bcd_in2=01000100 cout=1 sum=00000111
* bcd_in1=01100011 bcd_in2=01000101 cout=1 sum=00001000
* bcd_in1=01100011 bcd_in2=01000110 cout=1 sum=00001001
* bcd_in1=01100011 bcd_in2=01000111 cout=1 sum=00010000
* bcd_in1=01100011 bcd_in2=01001000 cout=1 sum=00010001
* bcd_in1=01100011 bcd_in2=01001001 cout=1 sum=00010010
* bcd_in1=01100011 bcd_in2=01010000 cout=1 sum=00010011
* bcd_in1=01100011 bcd_in2=01010001 cout=1 sum=00010100
* bcd_in1=01100011 bcd_in2=01010010 cout=1 sum=00010101
* bcd_in1=01100011 bcd_in2=01010011 cout=1 sum=00010110
* bcd_in1=01100011 bcd_in2=01010100 cout=1 sum=00010111
* bcd_in1=01100011 bcd_in2=01010101 cout=1 sum=00011000
* bcd_in1=01100011 bcd_in2=01010110 cout=1 sum=00011001
* bcd_in1=01100011 bcd_in2=01010111 cout=1 sum=00100000
* bcd_in1=01100011 bcd_in2=01011000 cout=1 sum=00100001
* bcd_in1=01100011 bcd_in2=01011001 cout=1 sum=00100010
* bcd_in1=01100011 bcd_in2=01100000 cout=1 sum=00100011
* bcd_in1=01100011 bcd_in2=01100001 cout=1 sum=00100100
* bcd_in1=01100011 bcd_in2=01100010 cout=1 sum=00100101
* bcd_in1=01100011 bcd_in2=01100011 cout=1 sum=00100110
* bcd_in1=01100011 bcd_in2=01100100 cout=1 sum=00100111
* bcd_in1=01100011 bcd_in2=01100101 cout=1 sum=00101000
* bcd_in1=01100011 bcd_in2=01100110 cout=1 sum=00101001
* bcd_in1=01100011 bcd_in2=01100111 cout=1 sum=00110000
* bcd_in1=01100011 bcd_in2=01101000 cout=1 sum=00110001
* bcd_in1=01100011 bcd_in2=01101001 cout=1 sum=00110010
* bcd_in1=01100011 bcd_in2=01110000 cout=1 sum=00110011
* bcd_in1=01100011 bcd_in2=01110001 cout=1 sum=00110100
* bcd_in1=01100011 bcd_in2=01110010 cout=1 sum=00110101
* bcd_in1=01100011 bcd_in2=01110011 cout=1 sum=00110110
* bcd_in1=01100011 bcd_in2=01110100 cout=1 sum=00110111
* bcd_in1=01100011 bcd_in2=01110101 cout=1 sum=00111000
* bcd_in1=01100011 bcd_in2=01110110 cout=1 sum=00111001
* bcd_in1=01100011 bcd_in2=01110111 cout=1 sum=01000000
* bcd_in1=01100011 bcd_in2=01111000 cout=1 sum=01000001
* bcd_in1=01100011 bcd_in2=01111001 cout=1 sum=01000010
* bcd_in1=01100011 bcd_in2=10000000 cout=1 sum=01000011
* bcd_in1=01100011 bcd_in2=10000001 cout=1 sum=01000100
* bcd_in1=01100011 bcd_in2=10000010 cout=1 sum=01000101
* bcd_in1=01100011 bcd_in2=10000011 cout=1 sum=01000110
* bcd_in1=01100011 bcd_in2=10000100 cout=1 sum=01000111
* bcd_in1=01100011 bcd_in2=10000101 cout=1 sum=01001000
* bcd_in1=01100011 bcd_in2=10000110 cout=1 sum=01001001
* bcd_in1=01100011 bcd_in2=10000111 cout=1 sum=01010000
* bcd_in1=01100011 bcd_in2=10001000 cout=1 sum=01010001
* bcd_in1=01100011 bcd_in2=10001001 cout=1 sum=01010010
* bcd_in1=01100011 bcd_in2=10010000 cout=1 sum=01010011
* bcd_in1=01100011 bcd_in2=10010001 cout=1 sum=01010100
* bcd_in1=01100011 bcd_in2=10010010 cout=1 sum=01010101
* bcd_in1=01100011 bcd_in2=10010011 cout=1 sum=01010110
* bcd_in1=01100011 bcd_in2=10010100 cout=1 sum=01010111
* bcd_in1=01100011 bcd_in2=10010101 cout=1 sum=01011000
* bcd_in1=01100011 bcd_in2=10010110 cout=1 sum=01011001
* bcd_in1=01100011 bcd_in2=10010111 cout=1 sum=01100000
* bcd_in1=01100011 bcd_in2=10011000 cout=1 sum=01100001
* bcd_in1=01100011 bcd_in2=10011001 cout=1 sum=01100010
* bcd_in1=01100100 bcd_in2=00000000 cout=0 sum=01100100
* bcd_in1=01100100 bcd_in2=00000001 cout=0 sum=01100101
* bcd_in1=01100100 bcd_in2=00000010 cout=0 sum=01100110
* bcd_in1=01100100 bcd_in2=00000011 cout=0 sum=01100111
* bcd_in1=01100100 bcd_in2=00000100 cout=0 sum=01101000
* bcd_in1=01100100 bcd_in2=00000101 cout=0 sum=01101001
* bcd_in1=01100100 bcd_in2=00000110 cout=0 sum=01110000
* bcd_in1=01100100 bcd_in2=00000111 cout=0 sum=01110001
* bcd_in1=01100100 bcd_in2=00001000 cout=0 sum=01110010
* bcd_in1=01100100 bcd_in2=00001001 cout=0 sum=01110011
* bcd_in1=01100100 bcd_in2=00010000 cout=0 sum=01110100
* bcd_in1=01100100 bcd_in2=00010001 cout=0 sum=01110101
* bcd_in1=01100100 bcd_in2=00010010 cout=0 sum=01110110
* bcd_in1=01100100 bcd_in2=00010011 cout=0 sum=01110111
* bcd_in1=01100100 bcd_in2=00010100 cout=0 sum=01111000
* bcd_in1=01100100 bcd_in2=00010101 cout=0 sum=01111001
* bcd_in1=01100100 bcd_in2=00010110 cout=0 sum=10000000
* bcd_in1=01100100 bcd_in2=00010111 cout=0 sum=10000001
* bcd_in1=01100100 bcd_in2=00011000 cout=0 sum=10000010
* bcd_in1=01100100 bcd_in2=00011001 cout=0 sum=10000011
* bcd_in1=01100100 bcd_in2=00100000 cout=0 sum=10000100
* bcd_in1=01100100 bcd_in2=00100001 cout=0 sum=10000101
* bcd_in1=01100100 bcd_in2=00100010 cout=0 sum=10000110
* bcd_in1=01100100 bcd_in2=00100011 cout=0 sum=10000111
* bcd_in1=01100100 bcd_in2=00100100 cout=0 sum=10001000
* bcd_in1=01100100 bcd_in2=00100101 cout=0 sum=10001001
* bcd_in1=01100100 bcd_in2=00100110 cout=0 sum=10010000
* bcd_in1=01100100 bcd_in2=00100111 cout=0 sum=10010001
* bcd_in1=01100100 bcd_in2=00101000 cout=0 sum=10010010
* bcd_in1=01100100 bcd_in2=00101001 cout=0 sum=10010011
* bcd_in1=01100100 bcd_in2=00110000 cout=0 sum=10010100
* bcd_in1=01100100 bcd_in2=00110001 cout=0 sum=10010101
* bcd_in1=01100100 bcd_in2=00110010 cout=0 sum=10010110
* bcd_in1=01100100 bcd_in2=00110011 cout=0 sum=10010111
* bcd_in1=01100100 bcd_in2=00110100 cout=0 sum=10011000
* bcd_in1=01100100 bcd_in2=00110101 cout=0 sum=10011001
* bcd_in1=01100100 bcd_in2=00110110 cout=1 sum=00000000
* bcd_in1=01100100 bcd_in2=00110111 cout=1 sum=00000001
* bcd_in1=01100100 bcd_in2=00111000 cout=1 sum=00000010
* bcd_in1=01100100 bcd_in2=00111001 cout=1 sum=00000011
* bcd_in1=01100100 bcd_in2=01000000 cout=1 sum=00000100
* bcd_in1=01100100 bcd_in2=01000001 cout=1 sum=00000101
* bcd_in1=01100100 bcd_in2=01000010 cout=1 sum=00000110
* bcd_in1=01100100 bcd_in2=01000011 cout=1 sum=00000111
* bcd_in1=01100100 bcd_in2=01000100 cout=1 sum=00001000
* bcd_in1=01100100 bcd_in2=01000101 cout=1 sum=00001001
* bcd_in1=01100100 bcd_in2=01000110 cout=1 sum=00010000
* bcd_in1=01100100 bcd_in2=01000111 cout=1 sum=00010001
* bcd_in1=01100100 bcd_in2=01001000 cout=1 sum=00010010
* bcd_in1=01100100 bcd_in2=01001001 cout=1 sum=00010011
* bcd_in1=01100100 bcd_in2=01010000 cout=1 sum=00010100
* bcd_in1=01100100 bcd_in2=01010001 cout=1 sum=00010101
* bcd_in1=01100100 bcd_in2=01010010 cout=1 sum=00010110
* bcd_in1=01100100 bcd_in2=01010011 cout=1 sum=00010111
* bcd_in1=01100100 bcd_in2=01010100 cout=1 sum=00011000
* bcd_in1=01100100 bcd_in2=01010101 cout=1 sum=00011001
* bcd_in1=01100100 bcd_in2=01010110 cout=1 sum=00100000
* bcd_in1=01100100 bcd_in2=01010111 cout=1 sum=00100001
* bcd_in1=01100100 bcd_in2=01011000 cout=1 sum=00100010
* bcd_in1=01100100 bcd_in2=01011001 cout=1 sum=00100011
* bcd_in1=01100100 bcd_in2=01100000 cout=1 sum=00100100
* bcd_in1=01100100 bcd_in2=01100001 cout=1 sum=00100101
* bcd_in1=01100100 bcd_in2=01100010 cout=1 sum=00100110
* bcd_in1=01100100 bcd_in2=01100011 cout=1 sum=00100111
* bcd_in1=01100100 bcd_in2=01100100 cout=1 sum=00101000
* bcd_in1=01100100 bcd_in2=01100101 cout=1 sum=00101001
* bcd_in1=01100100 bcd_in2=01100110 cout=1 sum=00110000
* bcd_in1=01100100 bcd_in2=01100111 cout=1 sum=00110001
* bcd_in1=01100100 bcd_in2=01101000 cout=1 sum=00110010
* bcd_in1=01100100 bcd_in2=01101001 cout=1 sum=00110011
* bcd_in1=01100100 bcd_in2=01110000 cout=1 sum=00110100
* bcd_in1=01100100 bcd_in2=01110001 cout=1 sum=00110101
* bcd_in1=01100100 bcd_in2=01110010 cout=1 sum=00110110
* bcd_in1=01100100 bcd_in2=01110011 cout=1 sum=00110111
* bcd_in1=01100100 bcd_in2=01110100 cout=1 sum=00111000
* bcd_in1=01100100 bcd_in2=01110101 cout=1 sum=00111001
* bcd_in1=01100100 bcd_in2=01110110 cout=1 sum=01000000
* bcd_in1=01100100 bcd_in2=01110111 cout=1 sum=01000001
* bcd_in1=01100100 bcd_in2=01111000 cout=1 sum=01000010
* bcd_in1=01100100 bcd_in2=01111001 cout=1 sum=01000011
* bcd_in1=01100100 bcd_in2=10000000 cout=1 sum=01000100
* bcd_in1=01100100 bcd_in2=10000001 cout=1 sum=01000101
* bcd_in1=01100100 bcd_in2=10000010 cout=1 sum=01000110
* bcd_in1=01100100 bcd_in2=10000011 cout=1 sum=01000111
* bcd_in1=01100100 bcd_in2=10000100 cout=1 sum=01001000
* bcd_in1=01100100 bcd_in2=10000101 cout=1 sum=01001001
* bcd_in1=01100100 bcd_in2=10000110 cout=1 sum=01010000
* bcd_in1=01100100 bcd_in2=10000111 cout=1 sum=01010001
* bcd_in1=01100100 bcd_in2=10001000 cout=1 sum=01010010
* bcd_in1=01100100 bcd_in2=10001001 cout=1 sum=01010011
* bcd_in1=01100100 bcd_in2=10010000 cout=1 sum=01010100
* bcd_in1=01100100 bcd_in2=10010001 cout=1 sum=01010101
* bcd_in1=01100100 bcd_in2=10010010 cout=1 sum=01010110
* bcd_in1=01100100 bcd_in2=10010011 cout=1 sum=01010111
* bcd_in1=01100100 bcd_in2=10010100 cout=1 sum=01011000
* bcd_in1=01100100 bcd_in2=10010101 cout=1 sum=01011001
* bcd_in1=01100100 bcd_in2=10010110 cout=1 sum=01100000
* bcd_in1=01100100 bcd_in2=10010111 cout=1 sum=01100001
* bcd_in1=01100100 bcd_in2=10011000 cout=1 sum=01100010
* bcd_in1=01100100 bcd_in2=10011001 cout=1 sum=01100011
* bcd_in1=01100101 bcd_in2=00000000 cout=0 sum=01100101
* bcd_in1=01100101 bcd_in2=00000001 cout=0 sum=01100110
* bcd_in1=01100101 bcd_in2=00000010 cout=0 sum=01100111
* bcd_in1=01100101 bcd_in2=00000011 cout=0 sum=01101000
* bcd_in1=01100101 bcd_in2=00000100 cout=0 sum=01101001
* bcd_in1=01100101 bcd_in2=00000101 cout=0 sum=01110000
* bcd_in1=01100101 bcd_in2=00000110 cout=0 sum=01110001
* bcd_in1=01100101 bcd_in2=00000111 cout=0 sum=01110010
* bcd_in1=01100101 bcd_in2=00001000 cout=0 sum=01110011
* bcd_in1=01100101 bcd_in2=00001001 cout=0 sum=01110100
* bcd_in1=01100101 bcd_in2=00010000 cout=0 sum=01110101
* bcd_in1=01100101 bcd_in2=00010001 cout=0 sum=01110110
* bcd_in1=01100101 bcd_in2=00010010 cout=0 sum=01110111
* bcd_in1=01100101 bcd_in2=00010011 cout=0 sum=01111000
* bcd_in1=01100101 bcd_in2=00010100 cout=0 sum=01111001
* bcd_in1=01100101 bcd_in2=00010101 cout=0 sum=10000000
* bcd_in1=01100101 bcd_in2=00010110 cout=0 sum=10000001
* bcd_in1=01100101 bcd_in2=00010111 cout=0 sum=10000010
* bcd_in1=01100101 bcd_in2=00011000 cout=0 sum=10000011
* bcd_in1=01100101 bcd_in2=00011001 cout=0 sum=10000100
* bcd_in1=01100101 bcd_in2=00100000 cout=0 sum=10000101
* bcd_in1=01100101 bcd_in2=00100001 cout=0 sum=10000110
* bcd_in1=01100101 bcd_in2=00100010 cout=0 sum=10000111
* bcd_in1=01100101 bcd_in2=00100011 cout=0 sum=10001000
* bcd_in1=01100101 bcd_in2=00100100 cout=0 sum=10001001
* bcd_in1=01100101 bcd_in2=00100101 cout=0 sum=10010000
* bcd_in1=01100101 bcd_in2=00100110 cout=0 sum=10010001
* bcd_in1=01100101 bcd_in2=00100111 cout=0 sum=10010010
* bcd_in1=01100101 bcd_in2=00101000 cout=0 sum=10010011
* bcd_in1=01100101 bcd_in2=00101001 cout=0 sum=10010100
* bcd_in1=01100101 bcd_in2=00110000 cout=0 sum=10010101
* bcd_in1=01100101 bcd_in2=00110001 cout=0 sum=10010110
* bcd_in1=01100101 bcd_in2=00110010 cout=0 sum=10010111
* bcd_in1=01100101 bcd_in2=00110011 cout=0 sum=10011000
* bcd_in1=01100101 bcd_in2=00110100 cout=0 sum=10011001
* bcd_in1=01100101 bcd_in2=00110101 cout=1 sum=00000000
* bcd_in1=01100101 bcd_in2=00110110 cout=1 sum=00000001
* bcd_in1=01100101 bcd_in2=00110111 cout=1 sum=00000010
* bcd_in1=01100101 bcd_in2=00111000 cout=1 sum=00000011
* bcd_in1=01100101 bcd_in2=00111001 cout=1 sum=00000100
* bcd_in1=01100101 bcd_in2=01000000 cout=1 sum=00000101
* bcd_in1=01100101 bcd_in2=01000001 cout=1 sum=00000110
* bcd_in1=01100101 bcd_in2=01000010 cout=1 sum=00000111
* bcd_in1=01100101 bcd_in2=01000011 cout=1 sum=00001000
* bcd_in1=01100101 bcd_in2=01000100 cout=1 sum=00001001
* bcd_in1=01100101 bcd_in2=01000101 cout=1 sum=00010000
* bcd_in1=01100101 bcd_in2=01000110 cout=1 sum=00010001
* bcd_in1=01100101 bcd_in2=01000111 cout=1 sum=00010010
* bcd_in1=01100101 bcd_in2=01001000 cout=1 sum=00010011
* bcd_in1=01100101 bcd_in2=01001001 cout=1 sum=00010100
* bcd_in1=01100101 bcd_in2=01010000 cout=1 sum=00010101
* bcd_in1=01100101 bcd_in2=01010001 cout=1 sum=00010110
* bcd_in1=01100101 bcd_in2=01010010 cout=1 sum=00010111
* bcd_in1=01100101 bcd_in2=01010011 cout=1 sum=00011000
* bcd_in1=01100101 bcd_in2=01010100 cout=1 sum=00011001
* bcd_in1=01100101 bcd_in2=01010101 cout=1 sum=00100000
* bcd_in1=01100101 bcd_in2=01010110 cout=1 sum=00100001
* bcd_in1=01100101 bcd_in2=01010111 cout=1 sum=00100010
* bcd_in1=01100101 bcd_in2=01011000 cout=1 sum=00100011
* bcd_in1=01100101 bcd_in2=01011001 cout=1 sum=00100100
* bcd_in1=01100101 bcd_in2=01100000 cout=1 sum=00100101
* bcd_in1=01100101 bcd_in2=01100001 cout=1 sum=00100110
* bcd_in1=01100101 bcd_in2=01100010 cout=1 sum=00100111
* bcd_in1=01100101 bcd_in2=01100011 cout=1 sum=00101000
* bcd_in1=01100101 bcd_in2=01100100 cout=1 sum=00101001
* bcd_in1=01100101 bcd_in2=01100101 cout=1 sum=00110000
* bcd_in1=01100101 bcd_in2=01100110 cout=1 sum=00110001
* bcd_in1=01100101 bcd_in2=01100111 cout=1 sum=00110010
* bcd_in1=01100101 bcd_in2=01101000 cout=1 sum=00110011
* bcd_in1=01100101 bcd_in2=01101001 cout=1 sum=00110100
* bcd_in1=01100101 bcd_in2=01110000 cout=1 sum=00110101
* bcd_in1=01100101 bcd_in2=01110001 cout=1 sum=00110110
* bcd_in1=01100101 bcd_in2=01110010 cout=1 sum=00110111
* bcd_in1=01100101 bcd_in2=01110011 cout=1 sum=00111000
* bcd_in1=01100101 bcd_in2=01110100 cout=1 sum=00111001
* bcd_in1=01100101 bcd_in2=01110101 cout=1 sum=01000000
* bcd_in1=01100101 bcd_in2=01110110 cout=1 sum=01000001
* bcd_in1=01100101 bcd_in2=01110111 cout=1 sum=01000010
* bcd_in1=01100101 bcd_in2=01111000 cout=1 sum=01000011
* bcd_in1=01100101 bcd_in2=01111001 cout=1 sum=01000100
* bcd_in1=01100101 bcd_in2=10000000 cout=1 sum=01000101
* bcd_in1=01100101 bcd_in2=10000001 cout=1 sum=01000110
* bcd_in1=01100101 bcd_in2=10000010 cout=1 sum=01000111
* bcd_in1=01100101 bcd_in2=10000011 cout=1 sum=01001000
* bcd_in1=01100101 bcd_in2=10000100 cout=1 sum=01001001
* bcd_in1=01100101 bcd_in2=10000101 cout=1 sum=01010000
* bcd_in1=01100101 bcd_in2=10000110 cout=1 sum=01010001
* bcd_in1=01100101 bcd_in2=10000111 cout=1 sum=01010010
* bcd_in1=01100101 bcd_in2=10001000 cout=1 sum=01010011
* bcd_in1=01100101 bcd_in2=10001001 cout=1 sum=01010100
* bcd_in1=01100101 bcd_in2=10010000 cout=1 sum=01010101
* bcd_in1=01100101 bcd_in2=10010001 cout=1 sum=01010110
* bcd_in1=01100101 bcd_in2=10010010 cout=1 sum=01010111
* bcd_in1=01100101 bcd_in2=10010011 cout=1 sum=01011000
* bcd_in1=01100101 bcd_in2=10010100 cout=1 sum=01011001
* bcd_in1=01100101 bcd_in2=10010101 cout=1 sum=01100000
* bcd_in1=01100101 bcd_in2=10010110 cout=1 sum=01100001
* bcd_in1=01100101 bcd_in2=10010111 cout=1 sum=01100010
* bcd_in1=01100101 bcd_in2=10011000 cout=1 sum=01100011
* bcd_in1=01100101 bcd_in2=10011001 cout=1 sum=01100100
* bcd_in1=01100110 bcd_in2=00000000 cout=0 sum=01100110
* bcd_in1=01100110 bcd_in2=00000001 cout=0 sum=01100111
* bcd_in1=01100110 bcd_in2=00000010 cout=0 sum=01101000
* bcd_in1=01100110 bcd_in2=00000011 cout=0 sum=01101001
* bcd_in1=01100110 bcd_in2=00000100 cout=0 sum=01110000
* bcd_in1=01100110 bcd_in2=00000101 cout=0 sum=01110001
* bcd_in1=01100110 bcd_in2=00000110 cout=0 sum=01110010
* bcd_in1=01100110 bcd_in2=00000111 cout=0 sum=01110011
* bcd_in1=01100110 bcd_in2=00001000 cout=0 sum=01110100
* bcd_in1=01100110 bcd_in2=00001001 cout=0 sum=01110101
* bcd_in1=01100110 bcd_in2=00010000 cout=0 sum=01110110
* bcd_in1=01100110 bcd_in2=00010001 cout=0 sum=01110111
* bcd_in1=01100110 bcd_in2=00010010 cout=0 sum=01111000
* bcd_in1=01100110 bcd_in2=00010011 cout=0 sum=01111001
* bcd_in1=01100110 bcd_in2=00010100 cout=0 sum=10000000
* bcd_in1=01100110 bcd_in2=00010101 cout=0 sum=10000001
* bcd_in1=01100110 bcd_in2=00010110 cout=0 sum=10000010
* bcd_in1=01100110 bcd_in2=00010111 cout=0 sum=10000011
* bcd_in1=01100110 bcd_in2=00011000 cout=0 sum=10000100
* bcd_in1=01100110 bcd_in2=00011001 cout=0 sum=10000101
* bcd_in1=01100110 bcd_in2=00100000 cout=0 sum=10000110
* bcd_in1=01100110 bcd_in2=00100001 cout=0 sum=10000111
* bcd_in1=01100110 bcd_in2=00100010 cout=0 sum=10001000
* bcd_in1=01100110 bcd_in2=00100011 cout=0 sum=10001001
* bcd_in1=01100110 bcd_in2=00100100 cout=0 sum=10010000
* bcd_in1=01100110 bcd_in2=00100101 cout=0 sum=10010001
* bcd_in1=01100110 bcd_in2=00100110 cout=0 sum=10010010
* bcd_in1=01100110 bcd_in2=00100111 cout=0 sum=10010011
* bcd_in1=01100110 bcd_in2=00101000 cout=0 sum=10010100
* bcd_in1=01100110 bcd_in2=00101001 cout=0 sum=10010101
* bcd_in1=01100110 bcd_in2=00110000 cout=0 sum=10010110
* bcd_in1=01100110 bcd_in2=00110001 cout=0 sum=10010111
* bcd_in1=01100110 bcd_in2=00110010 cout=0 sum=10011000
* bcd_in1=01100110 bcd_in2=00110011 cout=0 sum=10011001
* bcd_in1=01100110 bcd_in2=00110100 cout=1 sum=00000000
* bcd_in1=01100110 bcd_in2=00110101 cout=1 sum=00000001
* bcd_in1=01100110 bcd_in2=00110110 cout=1 sum=00000010
* bcd_in1=01100110 bcd_in2=00110111 cout=1 sum=00000011
* bcd_in1=01100110 bcd_in2=00111000 cout=1 sum=00000100
* bcd_in1=01100110 bcd_in2=00111001 cout=1 sum=00000101
* bcd_in1=01100110 bcd_in2=01000000 cout=1 sum=00000110
* bcd_in1=01100110 bcd_in2=01000001 cout=1 sum=00000111
* bcd_in1=01100110 bcd_in2=01000010 cout=1 sum=00001000
* bcd_in1=01100110 bcd_in2=01000011 cout=1 sum=00001001
* bcd_in1=01100110 bcd_in2=01000100 cout=1 sum=00010000
* bcd_in1=01100110 bcd_in2=01000101 cout=1 sum=00010001
* bcd_in1=01100110 bcd_in2=01000110 cout=1 sum=00010010
* bcd_in1=01100110 bcd_in2=01000111 cout=1 sum=00010011
* bcd_in1=01100110 bcd_in2=01001000 cout=1 sum=00010100
* bcd_in1=01100110 bcd_in2=01001001 cout=1 sum=00010101
* bcd_in1=01100110 bcd_in2=01010000 cout=1 sum=00010110
* bcd_in1=01100110 bcd_in2=01010001 cout=1 sum=00010111
* bcd_in1=01100110 bcd_in2=01010010 cout=1 sum=00011000
* bcd_in1=01100110 bcd_in2=01010011 cout=1 sum=00011001
* bcd_in1=01100110 bcd_in2=01010100 cout=1 sum=00100000
* bcd_in1=01100110 bcd_in2=01010101 cout=1 sum=00100001
* bcd_in1=01100110 bcd_in2=01010110 cout=1 sum=00100010
* bcd_in1=01100110 bcd_in2=01010111 cout=1 sum=00100011
* bcd_in1=01100110 bcd_in2=01011000 cout=1 sum=00100100
* bcd_in1=01100110 bcd_in2=01011001 cout=1 sum=00100101
* bcd_in1=01100110 bcd_in2=01100000 cout=1 sum=00100110
* bcd_in1=01100110 bcd_in2=01100001 cout=1 sum=00100111
* bcd_in1=01100110 bcd_in2=01100010 cout=1 sum=00101000
* bcd_in1=01100110 bcd_in2=01100011 cout=1 sum=00101001
* bcd_in1=01100110 bcd_in2=01100100 cout=1 sum=00110000
* bcd_in1=01100110 bcd_in2=01100101 cout=1 sum=00110001
* bcd_in1=01100110 bcd_in2=01100110 cout=1 sum=00110010
* bcd_in1=01100110 bcd_in2=01100111 cout=1 sum=00110011
* bcd_in1=01100110 bcd_in2=01101000 cout=1 sum=00110100
* bcd_in1=01100110 bcd_in2=01101001 cout=1 sum=00110101
* bcd_in1=01100110 bcd_in2=01110000 cout=1 sum=00110110
* bcd_in1=01100110 bcd_in2=01110001 cout=1 sum=00110111
* bcd_in1=01100110 bcd_in2=01110010 cout=1 sum=00111000
* bcd_in1=01100110 bcd_in2=01110011 cout=1 sum=00111001
* bcd_in1=01100110 bcd_in2=01110100 cout=1 sum=01000000
* bcd_in1=01100110 bcd_in2=01110101 cout=1 sum=01000001
* bcd_in1=01100110 bcd_in2=01110110 cout=1 sum=01000010
* bcd_in1=01100110 bcd_in2=01110111 cout=1 sum=01000011
* bcd_in1=01100110 bcd_in2=01111000 cout=1 sum=01000100
* bcd_in1=01100110 bcd_in2=01111001 cout=1 sum=01000101
* bcd_in1=01100110 bcd_in2=10000000 cout=1 sum=01000110
* bcd_in1=01100110 bcd_in2=10000001 cout=1 sum=01000111
* bcd_in1=01100110 bcd_in2=10000010 cout=1 sum=01001000
* bcd_in1=01100110 bcd_in2=10000011 cout=1 sum=01001001
* bcd_in1=01100110 bcd_in2=10000100 cout=1 sum=01010000
* bcd_in1=01100110 bcd_in2=10000101 cout=1 sum=01010001
* bcd_in1=01100110 bcd_in2=10000110 cout=1 sum=01010010
* bcd_in1=01100110 bcd_in2=10000111 cout=1 sum=01010011
* bcd_in1=01100110 bcd_in2=10001000 cout=1 sum=01010100
* bcd_in1=01100110 bcd_in2=10001001 cout=1 sum=01010101
* bcd_in1=01100110 bcd_in2=10010000 cout=1 sum=01010110
* bcd_in1=01100110 bcd_in2=10010001 cout=1 sum=01010111
* bcd_in1=01100110 bcd_in2=10010010 cout=1 sum=01011000
* bcd_in1=01100110 bcd_in2=10010011 cout=1 sum=01011001
* bcd_in1=01100110 bcd_in2=10010100 cout=1 sum=01100000
* bcd_in1=01100110 bcd_in2=10010101 cout=1 sum=01100001
* bcd_in1=01100110 bcd_in2=10010110 cout=1 sum=01100010
* bcd_in1=01100110 bcd_in2=10010111 cout=1 sum=01100011
* bcd_in1=01100110 bcd_in2=10011000 cout=1 sum=01100100
* bcd_in1=01100110 bcd_in2=10011001 cout=1 sum=01100101
* bcd_in1=01100111 bcd_in2=00000000 cout=0 sum=01100111
* bcd_in1=01100111 bcd_in2=00000001 cout=0 sum=01101000
* bcd_in1=01100111 bcd_in2=00000010 cout=0 sum=01101001
* bcd_in1=01100111 bcd_in2=00000011 cout=0 sum=01110000
* bcd_in1=01100111 bcd_in2=00000100 cout=0 sum=01110001
* bcd_in1=01100111 bcd_in2=00000101 cout=0 sum=01110010
* bcd_in1=01100111 bcd_in2=00000110 cout=0 sum=01110011
* bcd_in1=01100111 bcd_in2=00000111 cout=0 sum=01110100
* bcd_in1=01100111 bcd_in2=00001000 cout=0 sum=01110101
* bcd_in1=01100111 bcd_in2=00001001 cout=0 sum=01110110
* bcd_in1=01100111 bcd_in2=00010000 cout=0 sum=01110111
* bcd_in1=01100111 bcd_in2=00010001 cout=0 sum=01111000
* bcd_in1=01100111 bcd_in2=00010010 cout=0 sum=01111001
* bcd_in1=01100111 bcd_in2=00010011 cout=0 sum=10000000
* bcd_in1=01100111 bcd_in2=00010100 cout=0 sum=10000001
* bcd_in1=01100111 bcd_in2=00010101 cout=0 sum=10000010
* bcd_in1=01100111 bcd_in2=00010110 cout=0 sum=10000011
* bcd_in1=01100111 bcd_in2=00010111 cout=0 sum=10000100
* bcd_in1=01100111 bcd_in2=00011000 cout=0 sum=10000101
* bcd_in1=01100111 bcd_in2=00011001 cout=0 sum=10000110
* bcd_in1=01100111 bcd_in2=00100000 cout=0 sum=10000111
* bcd_in1=01100111 bcd_in2=00100001 cout=0 sum=10001000
* bcd_in1=01100111 bcd_in2=00100010 cout=0 sum=10001001
* bcd_in1=01100111 bcd_in2=00100011 cout=0 sum=10010000
* bcd_in1=01100111 bcd_in2=00100100 cout=0 sum=10010001
* bcd_in1=01100111 bcd_in2=00100101 cout=0 sum=10010010
* bcd_in1=01100111 bcd_in2=00100110 cout=0 sum=10010011
* bcd_in1=01100111 bcd_in2=00100111 cout=0 sum=10010100
* bcd_in1=01100111 bcd_in2=00101000 cout=0 sum=10010101
* bcd_in1=01100111 bcd_in2=00101001 cout=0 sum=10010110
* bcd_in1=01100111 bcd_in2=00110000 cout=0 sum=10010111
* bcd_in1=01100111 bcd_in2=00110001 cout=0 sum=10011000
* bcd_in1=01100111 bcd_in2=00110010 cout=0 sum=10011001
* bcd_in1=01100111 bcd_in2=00110011 cout=1 sum=00000000
* bcd_in1=01100111 bcd_in2=00110100 cout=1 sum=00000001
* bcd_in1=01100111 bcd_in2=00110101 cout=1 sum=00000010
* bcd_in1=01100111 bcd_in2=00110110 cout=1 sum=00000011
* bcd_in1=01100111 bcd_in2=00110111 cout=1 sum=00000100
* bcd_in1=01100111 bcd_in2=00111000 cout=1 sum=00000101
* bcd_in1=01100111 bcd_in2=00111001 cout=1 sum=00000110
* bcd_in1=01100111 bcd_in2=01000000 cout=1 sum=00000111
* bcd_in1=01100111 bcd_in2=01000001 cout=1 sum=00001000
* bcd_in1=01100111 bcd_in2=01000010 cout=1 sum=00001001
* bcd_in1=01100111 bcd_in2=01000011 cout=1 sum=00010000
* bcd_in1=01100111 bcd_in2=01000100 cout=1 sum=00010001
* bcd_in1=01100111 bcd_in2=01000101 cout=1 sum=00010010
* bcd_in1=01100111 bcd_in2=01000110 cout=1 sum=00010011
* bcd_in1=01100111 bcd_in2=01000111 cout=1 sum=00010100
* bcd_in1=01100111 bcd_in2=01001000 cout=1 sum=00010101
* bcd_in1=01100111 bcd_in2=01001001 cout=1 sum=00010110
* bcd_in1=01100111 bcd_in2=01010000 cout=1 sum=00010111
* bcd_in1=01100111 bcd_in2=01010001 cout=1 sum=00011000
* bcd_in1=01100111 bcd_in2=01010010 cout=1 sum=00011001
* bcd_in1=01100111 bcd_in2=01010011 cout=1 sum=00100000
* bcd_in1=01100111 bcd_in2=01010100 cout=1 sum=00100001
* bcd_in1=01100111 bcd_in2=01010101 cout=1 sum=00100010
* bcd_in1=01100111 bcd_in2=01010110 cout=1 sum=00100011
* bcd_in1=01100111 bcd_in2=01010111 cout=1 sum=00100100
* bcd_in1=01100111 bcd_in2=01011000 cout=1 sum=00100101
* bcd_in1=01100111 bcd_in2=01011001 cout=1 sum=00100110
* bcd_in1=01100111 bcd_in2=01100000 cout=1 sum=00100111
* bcd_in1=01100111 bcd_in2=01100001 cout=1 sum=00101000
* bcd_in1=01100111 bcd_in2=01100010 cout=1 sum=00101001
* bcd_in1=01100111 bcd_in2=01100011 cout=1 sum=00110000
* bcd_in1=01100111 bcd_in2=01100100 cout=1 sum=00110001
* bcd_in1=01100111 bcd_in2=01100101 cout=1 sum=00110010
* bcd_in1=01100111 bcd_in2=01100110 cout=1 sum=00110011
* bcd_in1=01100111 bcd_in2=01100111 cout=1 sum=00110100
* bcd_in1=01100111 bcd_in2=01101000 cout=1 sum=00110101
* bcd_in1=01100111 bcd_in2=01101001 cout=1 sum=00110110
* bcd_in1=01100111 bcd_in2=01110000 cout=1 sum=00110111
* bcd_in1=01100111 bcd_in2=01110001 cout=1 sum=00111000
* bcd_in1=01100111 bcd_in2=01110010 cout=1 sum=00111001
* bcd_in1=01100111 bcd_in2=01110011 cout=1 sum=01000000
* bcd_in1=01100111 bcd_in2=01110100 cout=1 sum=01000001
* bcd_in1=01100111 bcd_in2=01110101 cout=1 sum=01000010
* bcd_in1=01100111 bcd_in2=01110110 cout=1 sum=01000011
* bcd_in1=01100111 bcd_in2=01110111 cout=1 sum=01000100
* bcd_in1=01100111 bcd_in2=01111000 cout=1 sum=01000101
* bcd_in1=01100111 bcd_in2=01111001 cout=1 sum=01000110
* bcd_in1=01100111 bcd_in2=10000000 cout=1 sum=01000111
* bcd_in1=01100111 bcd_in2=10000001 cout=1 sum=01001000
* bcd_in1=01100111 bcd_in2=10000010 cout=1 sum=01001001
* bcd_in1=01100111 bcd_in2=10000011 cout=1 sum=01010000
* bcd_in1=01100111 bcd_in2=10000100 cout=1 sum=01010001
* bcd_in1=01100111 bcd_in2=10000101 cout=1 sum=01010010
* bcd_in1=01100111 bcd_in2=10000110 cout=1 sum=01010011
* bcd_in1=01100111 bcd_in2=10000111 cout=1 sum=01010100
* bcd_in1=01100111 bcd_in2=10001000 cout=1 sum=01010101
* bcd_in1=01100111 bcd_in2=10001001 cout=1 sum=01010110
* bcd_in1=01100111 bcd_in2=10010000 cout=1 sum=01010111
* bcd_in1=01100111 bcd_in2=10010001 cout=1 sum=01011000
* bcd_in1=01100111 bcd_in2=10010010 cout=1 sum=01011001
* bcd_in1=01100111 bcd_in2=10010011 cout=1 sum=01100000
* bcd_in1=01100111 bcd_in2=10010100 cout=1 sum=01100001
* bcd_in1=01100111 bcd_in2=10010101 cout=1 sum=01100010
* bcd_in1=01100111 bcd_in2=10010110 cout=1 sum=01100011
* bcd_in1=01100111 bcd_in2=10010111 cout=1 sum=01100100
* bcd_in1=01100111 bcd_in2=10011000 cout=1 sum=01100101
* bcd_in1=01100111 bcd_in2=10011001 cout=1 sum=01100110
* bcd_in1=01101000 bcd_in2=00000000 cout=0 sum=01101000
* bcd_in1=01101000 bcd_in2=00000001 cout=0 sum=01101001
* bcd_in1=01101000 bcd_in2=00000010 cout=0 sum=01110000
* bcd_in1=01101000 bcd_in2=00000011 cout=0 sum=01110001
* bcd_in1=01101000 bcd_in2=00000100 cout=0 sum=01110010
* bcd_in1=01101000 bcd_in2=00000101 cout=0 sum=01110011
* bcd_in1=01101000 bcd_in2=00000110 cout=0 sum=01110100
* bcd_in1=01101000 bcd_in2=00000111 cout=0 sum=01110101
* bcd_in1=01101000 bcd_in2=00001000 cout=0 sum=01110110
* bcd_in1=01101000 bcd_in2=00001001 cout=0 sum=01110111
* bcd_in1=01101000 bcd_in2=00010000 cout=0 sum=01111000
* bcd_in1=01101000 bcd_in2=00010001 cout=0 sum=01111001
* bcd_in1=01101000 bcd_in2=00010010 cout=0 sum=10000000
* bcd_in1=01101000 bcd_in2=00010011 cout=0 sum=10000001
* bcd_in1=01101000 bcd_in2=00010100 cout=0 sum=10000010
* bcd_in1=01101000 bcd_in2=00010101 cout=0 sum=10000011
* bcd_in1=01101000 bcd_in2=00010110 cout=0 sum=10000100
* bcd_in1=01101000 bcd_in2=00010111 cout=0 sum=10000101
* bcd_in1=01101000 bcd_in2=00011000 cout=0 sum=10000110
* bcd_in1=01101000 bcd_in2=00011001 cout=0 sum=10000111
* bcd_in1=01101000 bcd_in2=00100000 cout=0 sum=10001000
* bcd_in1=01101000 bcd_in2=00100001 cout=0 sum=10001001
* bcd_in1=01101000 bcd_in2=00100010 cout=0 sum=10010000
* bcd_in1=01101000 bcd_in2=00100011 cout=0 sum=10010001
* bcd_in1=01101000 bcd_in2=00100100 cout=0 sum=10010010
* bcd_in1=01101000 bcd_in2=00100101 cout=0 sum=10010011
* bcd_in1=01101000 bcd_in2=00100110 cout=0 sum=10010100
* bcd_in1=01101000 bcd_in2=00100111 cout=0 sum=10010101
* bcd_in1=01101000 bcd_in2=00101000 cout=0 sum=10010110
* bcd_in1=01101000 bcd_in2=00101001 cout=0 sum=10010111
* bcd_in1=01101000 bcd_in2=00110000 cout=0 sum=10011000
* bcd_in1=01101000 bcd_in2=00110001 cout=0 sum=10011001
* bcd_in1=01101000 bcd_in2=00110010 cout=1 sum=00000000
* bcd_in1=01101000 bcd_in2=00110011 cout=1 sum=00000001
* bcd_in1=01101000 bcd_in2=00110100 cout=1 sum=00000010
* bcd_in1=01101000 bcd_in2=00110101 cout=1 sum=00000011
* bcd_in1=01101000 bcd_in2=00110110 cout=1 sum=00000100
* bcd_in1=01101000 bcd_in2=00110111 cout=1 sum=00000101
* bcd_in1=01101000 bcd_in2=00111000 cout=1 sum=00000110
* bcd_in1=01101000 bcd_in2=00111001 cout=1 sum=00000111
* bcd_in1=01101000 bcd_in2=01000000 cout=1 sum=00001000
* bcd_in1=01101000 bcd_in2=01000001 cout=1 sum=00001001
* bcd_in1=01101000 bcd_in2=01000010 cout=1 sum=00010000
* bcd_in1=01101000 bcd_in2=01000011 cout=1 sum=00010001
* bcd_in1=01101000 bcd_in2=01000100 cout=1 sum=00010010
* bcd_in1=01101000 bcd_in2=01000101 cout=1 sum=00010011
* bcd_in1=01101000 bcd_in2=01000110 cout=1 sum=00010100
* bcd_in1=01101000 bcd_in2=01000111 cout=1 sum=00010101
* bcd_in1=01101000 bcd_in2=01001000 cout=1 sum=00010110
* bcd_in1=01101000 bcd_in2=01001001 cout=1 sum=00010111
* bcd_in1=01101000 bcd_in2=01010000 cout=1 sum=00011000
* bcd_in1=01101000 bcd_in2=01010001 cout=1 sum=00011001
* bcd_in1=01101000 bcd_in2=01010010 cout=1 sum=00100000
* bcd_in1=01101000 bcd_in2=01010011 cout=1 sum=00100001
* bcd_in1=01101000 bcd_in2=01010100 cout=1 sum=00100010
* bcd_in1=01101000 bcd_in2=01010101 cout=1 sum=00100011
* bcd_in1=01101000 bcd_in2=01010110 cout=1 sum=00100100
* bcd_in1=01101000 bcd_in2=01010111 cout=1 sum=00100101
* bcd_in1=01101000 bcd_in2=01011000 cout=1 sum=00100110
* bcd_in1=01101000 bcd_in2=01011001 cout=1 sum=00100111
* bcd_in1=01101000 bcd_in2=01100000 cout=1 sum=00101000
* bcd_in1=01101000 bcd_in2=01100001 cout=1 sum=00101001
* bcd_in1=01101000 bcd_in2=01100010 cout=1 sum=00110000
* bcd_in1=01101000 bcd_in2=01100011 cout=1 sum=00110001
* bcd_in1=01101000 bcd_in2=01100100 cout=1 sum=00110010
* bcd_in1=01101000 bcd_in2=01100101 cout=1 sum=00110011
* bcd_in1=01101000 bcd_in2=01100110 cout=1 sum=00110100
* bcd_in1=01101000 bcd_in2=01100111 cout=1 sum=00110101
* bcd_in1=01101000 bcd_in2=01101000 cout=1 sum=00110110
* bcd_in1=01101000 bcd_in2=01101001 cout=1 sum=00110111
* bcd_in1=01101000 bcd_in2=01110000 cout=1 sum=00111000
* bcd_in1=01101000 bcd_in2=01110001 cout=1 sum=00111001
* bcd_in1=01101000 bcd_in2=01110010 cout=1 sum=01000000
* bcd_in1=01101000 bcd_in2=01110011 cout=1 sum=01000001
* bcd_in1=01101000 bcd_in2=01110100 cout=1 sum=01000010
* bcd_in1=01101000 bcd_in2=01110101 cout=1 sum=01000011
* bcd_in1=01101000 bcd_in2=01110110 cout=1 sum=01000100
* bcd_in1=01101000 bcd_in2=01110111 cout=1 sum=01000101
* bcd_in1=01101000 bcd_in2=01111000 cout=1 sum=01000110
* bcd_in1=01101000 bcd_in2=01111001 cout=1 sum=01000111
* bcd_in1=01101000 bcd_in2=10000000 cout=1 sum=01001000
* bcd_in1=01101000 bcd_in2=10000001 cout=1 sum=01001001
* bcd_in1=01101000 bcd_in2=10000010 cout=1 sum=01010000
* bcd_in1=01101000 bcd_in2=10000011 cout=1 sum=01010001
* bcd_in1=01101000 bcd_in2=10000100 cout=1 sum=01010010
* bcd_in1=01101000 bcd_in2=10000101 cout=1 sum=01010011
* bcd_in1=01101000 bcd_in2=10000110 cout=1 sum=01010100
* bcd_in1=01101000 bcd_in2=10000111 cout=1 sum=01010101
* bcd_in1=01101000 bcd_in2=10001000 cout=1 sum=01010110
* bcd_in1=01101000 bcd_in2=10001001 cout=1 sum=01010111
* bcd_in1=01101000 bcd_in2=10010000 cout=1 sum=01011000
* bcd_in1=01101000 bcd_in2=10010001 cout=1 sum=01011001
* bcd_in1=01101000 bcd_in2=10010010 cout=1 sum=01100000
* bcd_in1=01101000 bcd_in2=10010011 cout=1 sum=01100001
* bcd_in1=01101000 bcd_in2=10010100 cout=1 sum=01100010
* bcd_in1=01101000 bcd_in2=10010101 cout=1 sum=01100011
* bcd_in1=01101000 bcd_in2=10010110 cout=1 sum=01100100
* bcd_in1=01101000 bcd_in2=10010111 cout=1 sum=01100101
* bcd_in1=01101000 bcd_in2=10011000 cout=1 sum=01100110
* bcd_in1=01101000 bcd_in2=10011001 cout=1 sum=01100111
* bcd_in1=01101001 bcd_in2=00000000 cout=0 sum=01101001
* bcd_in1=01101001 bcd_in2=00000001 cout=0 sum=01110000
* bcd_in1=01101001 bcd_in2=00000010 cout=0 sum=01110001
* bcd_in1=01101001 bcd_in2=00000011 cout=0 sum=01110010
* bcd_in1=01101001 bcd_in2=00000100 cout=0 sum=01110011
* bcd_in1=01101001 bcd_in2=00000101 cout=0 sum=01110100
* bcd_in1=01101001 bcd_in2=00000110 cout=0 sum=01110101
* bcd_in1=01101001 bcd_in2=00000111 cout=0 sum=01110110
* bcd_in1=01101001 bcd_in2=00001000 cout=0 sum=01110111
* bcd_in1=01101001 bcd_in2=00001001 cout=0 sum=01111000
* bcd_in1=01101001 bcd_in2=00010000 cout=0 sum=01111001
* bcd_in1=01101001 bcd_in2=00010001 cout=0 sum=10000000
* bcd_in1=01101001 bcd_in2=00010010 cout=0 sum=10000001
* bcd_in1=01101001 bcd_in2=00010011 cout=0 sum=10000010
* bcd_in1=01101001 bcd_in2=00010100 cout=0 sum=10000011
* bcd_in1=01101001 bcd_in2=00010101 cout=0 sum=10000100
* bcd_in1=01101001 bcd_in2=00010110 cout=0 sum=10000101
* bcd_in1=01101001 bcd_in2=00010111 cout=0 sum=10000110
* bcd_in1=01101001 bcd_in2=00011000 cout=0 sum=10000111
* bcd_in1=01101001 bcd_in2=00011001 cout=0 sum=10001000
* bcd_in1=01101001 bcd_in2=00100000 cout=0 sum=10001001
* bcd_in1=01101001 bcd_in2=00100001 cout=0 sum=10010000
* bcd_in1=01101001 bcd_in2=00100010 cout=0 sum=10010001
* bcd_in1=01101001 bcd_in2=00100011 cout=0 sum=10010010
* bcd_in1=01101001 bcd_in2=00100100 cout=0 sum=10010011
* bcd_in1=01101001 bcd_in2=00100101 cout=0 sum=10010100
* bcd_in1=01101001 bcd_in2=00100110 cout=0 sum=10010101
* bcd_in1=01101001 bcd_in2=00100111 cout=0 sum=10010110
* bcd_in1=01101001 bcd_in2=00101000 cout=0 sum=10010111
* bcd_in1=01101001 bcd_in2=00101001 cout=0 sum=10011000
* bcd_in1=01101001 bcd_in2=00110000 cout=0 sum=10011001
* bcd_in1=01101001 bcd_in2=00110001 cout=1 sum=00000000
* bcd_in1=01101001 bcd_in2=00110010 cout=1 sum=00000001
* bcd_in1=01101001 bcd_in2=00110011 cout=1 sum=00000010
* bcd_in1=01101001 bcd_in2=00110100 cout=1 sum=00000011
* bcd_in1=01101001 bcd_in2=00110101 cout=1 sum=00000100
* bcd_in1=01101001 bcd_in2=00110110 cout=1 sum=00000101
* bcd_in1=01101001 bcd_in2=00110111 cout=1 sum=00000110
* bcd_in1=01101001 bcd_in2=00111000 cout=1 sum=00000111
* bcd_in1=01101001 bcd_in2=00111001 cout=1 sum=00001000
* bcd_in1=01101001 bcd_in2=01000000 cout=1 sum=00001001
* bcd_in1=01101001 bcd_in2=01000001 cout=1 sum=00010000
* bcd_in1=01101001 bcd_in2=01000010 cout=1 sum=00010001
* bcd_in1=01101001 bcd_in2=01000011 cout=1 sum=00010010
* bcd_in1=01101001 bcd_in2=01000100 cout=1 sum=00010011
* bcd_in1=01101001 bcd_in2=01000101 cout=1 sum=00010100
* bcd_in1=01101001 bcd_in2=01000110 cout=1 sum=00010101
* bcd_in1=01101001 bcd_in2=01000111 cout=1 sum=00010110
* bcd_in1=01101001 bcd_in2=01001000 cout=1 sum=00010111
* bcd_in1=01101001 bcd_in2=01001001 cout=1 sum=00011000
* bcd_in1=01101001 bcd_in2=01010000 cout=1 sum=00011001
* bcd_in1=01101001 bcd_in2=01010001 cout=1 sum=00100000
* bcd_in1=01101001 bcd_in2=01010010 cout=1 sum=00100001
* bcd_in1=01101001 bcd_in2=01010011 cout=1 sum=00100010
* bcd_in1=01101001 bcd_in2=01010100 cout=1 sum=00100011
* bcd_in1=01101001 bcd_in2=01010101 cout=1 sum=00100100
* bcd_in1=01101001 bcd_in2=01010110 cout=1 sum=00100101
* bcd_in1=01101001 bcd_in2=01010111 cout=1 sum=00100110
* bcd_in1=01101001 bcd_in2=01011000 cout=1 sum=00100111
* bcd_in1=01101001 bcd_in2=01011001 cout=1 sum=00101000
* bcd_in1=01101001 bcd_in2=01100000 cout=1 sum=00101001
* bcd_in1=01101001 bcd_in2=01100001 cout=1 sum=00110000
* bcd_in1=01101001 bcd_in2=01100010 cout=1 sum=00110001
* bcd_in1=01101001 bcd_in2=01100011 cout=1 sum=00110010
* bcd_in1=01101001 bcd_in2=01100100 cout=1 sum=00110011
* bcd_in1=01101001 bcd_in2=01100101 cout=1 sum=00110100
* bcd_in1=01101001 bcd_in2=01100110 cout=1 sum=00110101
* bcd_in1=01101001 bcd_in2=01100111 cout=1 sum=00110110
* bcd_in1=01101001 bcd_in2=01101000 cout=1 sum=00110111
* bcd_in1=01101001 bcd_in2=01101001 cout=1 sum=00111000
* bcd_in1=01101001 bcd_in2=01110000 cout=1 sum=00111001
* bcd_in1=01101001 bcd_in2=01110001 cout=1 sum=01000000
* bcd_in1=01101001 bcd_in2=01110010 cout=1 sum=01000001
* bcd_in1=01101001 bcd_in2=01110011 cout=1 sum=01000010
* bcd_in1=01101001 bcd_in2=01110100 cout=1 sum=01000011
* bcd_in1=01101001 bcd_in2=01110101 cout=1 sum=01000100
* bcd_in1=01101001 bcd_in2=01110110 cout=1 sum=01000101
* bcd_in1=01101001 bcd_in2=01110111 cout=1 sum=01000110
* bcd_in1=01101001 bcd_in2=01111000 cout=1 sum=01000111
* bcd_in1=01101001 bcd_in2=01111001 cout=1 sum=01001000
* bcd_in1=01101001 bcd_in2=10000000 cout=1 sum=01001001
* bcd_in1=01101001 bcd_in2=10000001 cout=1 sum=01010000
* bcd_in1=01101001 bcd_in2=10000010 cout=1 sum=01010001
* bcd_in1=01101001 bcd_in2=10000011 cout=1 sum=01010010
* bcd_in1=01101001 bcd_in2=10000100 cout=1 sum=01010011
* bcd_in1=01101001 bcd_in2=10000101 cout=1 sum=01010100
* bcd_in1=01101001 bcd_in2=10000110 cout=1 sum=01010101
* bcd_in1=01101001 bcd_in2=10000111 cout=1 sum=01010110
* bcd_in1=01101001 bcd_in2=10001000 cout=1 sum=01010111
* bcd_in1=01101001 bcd_in2=10001001 cout=1 sum=01011000
* bcd_in1=01101001 bcd_in2=10010000 cout=1 sum=01011001
* bcd_in1=01101001 bcd_in2=10010001 cout=1 sum=01100000
* bcd_in1=01101001 bcd_in2=10010010 cout=1 sum=01100001
* bcd_in1=01101001 bcd_in2=10010011 cout=1 sum=01100010
* bcd_in1=01101001 bcd_in2=10010100 cout=1 sum=01100011
* bcd_in1=01101001 bcd_in2=10010101 cout=1 sum=01100100
* bcd_in1=01101001 bcd_in2=10010110 cout=1 sum=01100101
* bcd_in1=01101001 bcd_in2=10010111 cout=1 sum=01100110
* bcd_in1=01101001 bcd_in2=10011000 cout=1 sum=01100111
* bcd_in1=01101001 bcd_in2=10011001 cout=1 sum=01101000
* bcd_in1=01110000 bcd_in2=00000000 cout=0 sum=01110000
* bcd_in1=01110000 bcd_in2=00000001 cout=0 sum=01110001
* bcd_in1=01110000 bcd_in2=00000010 cout=0 sum=01110010
* bcd_in1=01110000 bcd_in2=00000011 cout=0 sum=01110011
* bcd_in1=01110000 bcd_in2=00000100 cout=0 sum=01110100
* bcd_in1=01110000 bcd_in2=00000101 cout=0 sum=01110101
* bcd_in1=01110000 bcd_in2=00000110 cout=0 sum=01110110
* bcd_in1=01110000 bcd_in2=00000111 cout=0 sum=01110111
* bcd_in1=01110000 bcd_in2=00001000 cout=0 sum=01111000
* bcd_in1=01110000 bcd_in2=00001001 cout=0 sum=01111001
* bcd_in1=01110000 bcd_in2=00010000 cout=0 sum=10000000
* bcd_in1=01110000 bcd_in2=00010001 cout=0 sum=10000001
* bcd_in1=01110000 bcd_in2=00010010 cout=0 sum=10000010
* bcd_in1=01110000 bcd_in2=00010011 cout=0 sum=10000011
* bcd_in1=01110000 bcd_in2=00010100 cout=0 sum=10000100
* bcd_in1=01110000 bcd_in2=00010101 cout=0 sum=10000101
* bcd_in1=01110000 bcd_in2=00010110 cout=0 sum=10000110
* bcd_in1=01110000 bcd_in2=00010111 cout=0 sum=10000111
* bcd_in1=01110000 bcd_in2=00011000 cout=0 sum=10001000
* bcd_in1=01110000 bcd_in2=00011001 cout=0 sum=10001001
* bcd_in1=01110000 bcd_in2=00100000 cout=0 sum=10010000
* bcd_in1=01110000 bcd_in2=00100001 cout=0 sum=10010001
* bcd_in1=01110000 bcd_in2=00100010 cout=0 sum=10010010
* bcd_in1=01110000 bcd_in2=00100011 cout=0 sum=10010011
* bcd_in1=01110000 bcd_in2=00100100 cout=0 sum=10010100
* bcd_in1=01110000 bcd_in2=00100101 cout=0 sum=10010101
* bcd_in1=01110000 bcd_in2=00100110 cout=0 sum=10010110
* bcd_in1=01110000 bcd_in2=00100111 cout=0 sum=10010111
* bcd_in1=01110000 bcd_in2=00101000 cout=0 sum=10011000
* bcd_in1=01110000 bcd_in2=00101001 cout=0 sum=10011001
* bcd_in1=01110000 bcd_in2=00110000 cout=1 sum=00000000
* bcd_in1=01110000 bcd_in2=00110001 cout=1 sum=00000001
* bcd_in1=01110000 bcd_in2=00110010 cout=1 sum=00000010
* bcd_in1=01110000 bcd_in2=00110011 cout=1 sum=00000011
* bcd_in1=01110000 bcd_in2=00110100 cout=1 sum=00000100
* bcd_in1=01110000 bcd_in2=00110101 cout=1 sum=00000101
* bcd_in1=01110000 bcd_in2=00110110 cout=1 sum=00000110
* bcd_in1=01110000 bcd_in2=00110111 cout=1 sum=00000111
* bcd_in1=01110000 bcd_in2=00111000 cout=1 sum=00001000
* bcd_in1=01110000 bcd_in2=00111001 cout=1 sum=00001001
* bcd_in1=01110000 bcd_in2=01000000 cout=1 sum=00010000
* bcd_in1=01110000 bcd_in2=01000001 cout=1 sum=00010001
* bcd_in1=01110000 bcd_in2=01000010 cout=1 sum=00010010
* bcd_in1=01110000 bcd_in2=01000011 cout=1 sum=00010011
* bcd_in1=01110000 bcd_in2=01000100 cout=1 sum=00010100
* bcd_in1=01110000 bcd_in2=01000101 cout=1 sum=00010101
* bcd_in1=01110000 bcd_in2=01000110 cout=1 sum=00010110
* bcd_in1=01110000 bcd_in2=01000111 cout=1 sum=00010111
* bcd_in1=01110000 bcd_in2=01001000 cout=1 sum=00011000
* bcd_in1=01110000 bcd_in2=01001001 cout=1 sum=00011001
* bcd_in1=01110000 bcd_in2=01010000 cout=1 sum=00100000
* bcd_in1=01110000 bcd_in2=01010001 cout=1 sum=00100001
* bcd_in1=01110000 bcd_in2=01010010 cout=1 sum=00100010
* bcd_in1=01110000 bcd_in2=01010011 cout=1 sum=00100011
* bcd_in1=01110000 bcd_in2=01010100 cout=1 sum=00100100
* bcd_in1=01110000 bcd_in2=01010101 cout=1 sum=00100101
* bcd_in1=01110000 bcd_in2=01010110 cout=1 sum=00100110
* bcd_in1=01110000 bcd_in2=01010111 cout=1 sum=00100111
* bcd_in1=01110000 bcd_in2=01011000 cout=1 sum=00101000
* bcd_in1=01110000 bcd_in2=01011001 cout=1 sum=00101001
* bcd_in1=01110000 bcd_in2=01100000 cout=1 sum=00110000
* bcd_in1=01110000 bcd_in2=01100001 cout=1 sum=00110001
* bcd_in1=01110000 bcd_in2=01100010 cout=1 sum=00110010
* bcd_in1=01110000 bcd_in2=01100011 cout=1 sum=00110011
* bcd_in1=01110000 bcd_in2=01100100 cout=1 sum=00110100
* bcd_in1=01110000 bcd_in2=01100101 cout=1 sum=00110101
* bcd_in1=01110000 bcd_in2=01100110 cout=1 sum=00110110
* bcd_in1=01110000 bcd_in2=01100111 cout=1 sum=00110111
* bcd_in1=01110000 bcd_in2=01101000 cout=1 sum=00111000
* bcd_in1=01110000 bcd_in2=01101001 cout=1 sum=00111001
* bcd_in1=01110000 bcd_in2=01110000 cout=1 sum=01000000
* bcd_in1=01110000 bcd_in2=01110001 cout=1 sum=01000001
* bcd_in1=01110000 bcd_in2=01110010 cout=1 sum=01000010
* bcd_in1=01110000 bcd_in2=01110011 cout=1 sum=01000011
* bcd_in1=01110000 bcd_in2=01110100 cout=1 sum=01000100
* bcd_in1=01110000 bcd_in2=01110101 cout=1 sum=01000101
* bcd_in1=01110000 bcd_in2=01110110 cout=1 sum=01000110
* bcd_in1=01110000 bcd_in2=01110111 cout=1 sum=01000111
* bcd_in1=01110000 bcd_in2=01111000 cout=1 sum=01001000
* bcd_in1=01110000 bcd_in2=01111001 cout=1 sum=01001001
* bcd_in1=01110000 bcd_in2=10000000 cout=1 sum=01010000
* bcd_in1=01110000 bcd_in2=10000001 cout=1 sum=01010001
* bcd_in1=01110000 bcd_in2=10000010 cout=1 sum=01010010
* bcd_in1=01110000 bcd_in2=10000011 cout=1 sum=01010011
* bcd_in1=01110000 bcd_in2=10000100 cout=1 sum=01010100
* bcd_in1=01110000 bcd_in2=10000101 cout=1 sum=01010101
* bcd_in1=01110000 bcd_in2=10000110 cout=1 sum=01010110
* bcd_in1=01110000 bcd_in2=10000111 cout=1 sum=01010111
* bcd_in1=01110000 bcd_in2=10001000 cout=1 sum=01011000
* bcd_in1=01110000 bcd_in2=10001001 cout=1 sum=01011001
* bcd_in1=01110000 bcd_in2=10010000 cout=1 sum=01100000
* bcd_in1=01110000 bcd_in2=10010001 cout=1 sum=01100001
* bcd_in1=01110000 bcd_in2=10010010 cout=1 sum=01100010
* bcd_in1=01110000 bcd_in2=10010011 cout=1 sum=01100011
* bcd_in1=01110000 bcd_in2=10010100 cout=1 sum=01100100
* bcd_in1=01110000 bcd_in2=10010101 cout=1 sum=01100101
* bcd_in1=01110000 bcd_in2=10010110 cout=1 sum=01100110
* bcd_in1=01110000 bcd_in2=10010111 cout=1 sum=01100111
* bcd_in1=01110000 bcd_in2=10011000 cout=1 sum=01101000
* bcd_in1=01110000 bcd_in2=10011001 cout=1 sum=01101001
* bcd_in1=01110001 bcd_in2=00000000 cout=0 sum=01110001
* bcd_in1=01110001 bcd_in2=00000001 cout=0 sum=01110010
* bcd_in1=01110001 bcd_in2=00000010 cout=0 sum=01110011
* bcd_in1=01110001 bcd_in2=00000011 cout=0 sum=01110100
* bcd_in1=01110001 bcd_in2=00000100 cout=0 sum=01110101
* bcd_in1=01110001 bcd_in2=00000101 cout=0 sum=01110110
* bcd_in1=01110001 bcd_in2=00000110 cout=0 sum=01110111
* bcd_in1=01110001 bcd_in2=00000111 cout=0 sum=01111000
* bcd_in1=01110001 bcd_in2=00001000 cout=0 sum=01111001
* bcd_in1=01110001 bcd_in2=00001001 cout=0 sum=10000000
* bcd_in1=01110001 bcd_in2=00010000 cout=0 sum=10000001
* bcd_in1=01110001 bcd_in2=00010001 cout=0 sum=10000010
* bcd_in1=01110001 bcd_in2=00010010 cout=0 sum=10000011
* bcd_in1=01110001 bcd_in2=00010011 cout=0 sum=10000100
* bcd_in1=01110001 bcd_in2=00010100 cout=0 sum=10000101
* bcd_in1=01110001 bcd_in2=00010101 cout=0 sum=10000110
* bcd_in1=01110001 bcd_in2=00010110 cout=0 sum=10000111
* bcd_in1=01110001 bcd_in2=00010111 cout=0 sum=10001000
* bcd_in1=01110001 bcd_in2=00011000 cout=0 sum=10001001
* bcd_in1=01110001 bcd_in2=00011001 cout=0 sum=10010000
* bcd_in1=01110001 bcd_in2=00100000 cout=0 sum=10010001
* bcd_in1=01110001 bcd_in2=00100001 cout=0 sum=10010010
* bcd_in1=01110001 bcd_in2=00100010 cout=0 sum=10010011
* bcd_in1=01110001 bcd_in2=00100011 cout=0 sum=10010100
* bcd_in1=01110001 bcd_in2=00100100 cout=0 sum=10010101
* bcd_in1=01110001 bcd_in2=00100101 cout=0 sum=10010110
* bcd_in1=01110001 bcd_in2=00100110 cout=0 sum=10010111
* bcd_in1=01110001 bcd_in2=00100111 cout=0 sum=10011000
* bcd_in1=01110001 bcd_in2=00101000 cout=0 sum=10011001
* bcd_in1=01110001 bcd_in2=00101001 cout=1 sum=00000000
* bcd_in1=01110001 bcd_in2=00110000 cout=1 sum=00000001
* bcd_in1=01110001 bcd_in2=00110001 cout=1 sum=00000010
* bcd_in1=01110001 bcd_in2=00110010 cout=1 sum=00000011
* bcd_in1=01110001 bcd_in2=00110011 cout=1 sum=00000100
* bcd_in1=01110001 bcd_in2=00110100 cout=1 sum=00000101
* bcd_in1=01110001 bcd_in2=00110101 cout=1 sum=00000110
* bcd_in1=01110001 bcd_in2=00110110 cout=1 sum=00000111
* bcd_in1=01110001 bcd_in2=00110111 cout=1 sum=00001000
* bcd_in1=01110001 bcd_in2=00111000 cout=1 sum=00001001
* bcd_in1=01110001 bcd_in2=00111001 cout=1 sum=00010000
* bcd_in1=01110001 bcd_in2=01000000 cout=1 sum=00010001
* bcd_in1=01110001 bcd_in2=01000001 cout=1 sum=00010010
* bcd_in1=01110001 bcd_in2=01000010 cout=1 sum=00010011
* bcd_in1=01110001 bcd_in2=01000011 cout=1 sum=00010100
* bcd_in1=01110001 bcd_in2=01000100 cout=1 sum=00010101
* bcd_in1=01110001 bcd_in2=01000101 cout=1 sum=00010110
* bcd_in1=01110001 bcd_in2=01000110 cout=1 sum=00010111
* bcd_in1=01110001 bcd_in2=01000111 cout=1 sum=00011000
* bcd_in1=01110001 bcd_in2=01001000 cout=1 sum=00011001
* bcd_in1=01110001 bcd_in2=01001001 cout=1 sum=00100000
* bcd_in1=01110001 bcd_in2=01010000 cout=1 sum=00100001
* bcd_in1=01110001 bcd_in2=01010001 cout=1 sum=00100010
* bcd_in1=01110001 bcd_in2=01010010 cout=1 sum=00100011
* bcd_in1=01110001 bcd_in2=01010011 cout=1 sum=00100100
* bcd_in1=01110001 bcd_in2=01010100 cout=1 sum=00100101
* bcd_in1=01110001 bcd_in2=01010101 cout=1 sum=00100110
* bcd_in1=01110001 bcd_in2=01010110 cout=1 sum=00100111
* bcd_in1=01110001 bcd_in2=01010111 cout=1 sum=00101000
* bcd_in1=01110001 bcd_in2=01011000 cout=1 sum=00101001
* bcd_in1=01110001 bcd_in2=01011001 cout=1 sum=00110000
* bcd_in1=01110001 bcd_in2=01100000 cout=1 sum=00110001
* bcd_in1=01110001 bcd_in2=01100001 cout=1 sum=00110010
* bcd_in1=01110001 bcd_in2=01100010 cout=1 sum=00110011
* bcd_in1=01110001 bcd_in2=01100011 cout=1 sum=00110100
* bcd_in1=01110001 bcd_in2=01100100 cout=1 sum=00110101
* bcd_in1=01110001 bcd_in2=01100101 cout=1 sum=00110110
* bcd_in1=01110001 bcd_in2=01100110 cout=1 sum=00110111
* bcd_in1=01110001 bcd_in2=01100111 cout=1 sum=00111000
* bcd_in1=01110001 bcd_in2=01101000 cout=1 sum=00111001
* bcd_in1=01110001 bcd_in2=01101001 cout=1 sum=01000000
* bcd_in1=01110001 bcd_in2=01110000 cout=1 sum=01000001
* bcd_in1=01110001 bcd_in2=01110001 cout=1 sum=01000010
* bcd_in1=01110001 bcd_in2=01110010 cout=1 sum=01000011
* bcd_in1=01110001 bcd_in2=01110011 cout=1 sum=01000100
* bcd_in1=01110001 bcd_in2=01110100 cout=1 sum=01000101
* bcd_in1=01110001 bcd_in2=01110101 cout=1 sum=01000110
* bcd_in1=01110001 bcd_in2=01110110 cout=1 sum=01000111
* bcd_in1=01110001 bcd_in2=01110111 cout=1 sum=01001000
* bcd_in1=01110001 bcd_in2=01111000 cout=1 sum=01001001
* bcd_in1=01110001 bcd_in2=01111001 cout=1 sum=01010000
* bcd_in1=01110001 bcd_in2=10000000 cout=1 sum=01010001
* bcd_in1=01110001 bcd_in2=10000001 cout=1 sum=01010010
* bcd_in1=01110001 bcd_in2=10000010 cout=1 sum=01010011
* bcd_in1=01110001 bcd_in2=10000011 cout=1 sum=01010100
* bcd_in1=01110001 bcd_in2=10000100 cout=1 sum=01010101
* bcd_in1=01110001 bcd_in2=10000101 cout=1 sum=01010110
* bcd_in1=01110001 bcd_in2=10000110 cout=1 sum=01010111
* bcd_in1=01110001 bcd_in2=10000111 cout=1 sum=01011000
* bcd_in1=01110001 bcd_in2=10001000 cout=1 sum=01011001
* bcd_in1=01110001 bcd_in2=10001001 cout=1 sum=01100000
* bcd_in1=01110001 bcd_in2=10010000 cout=1 sum=01100001
* bcd_in1=01110001 bcd_in2=10010001 cout=1 sum=01100010
* bcd_in1=01110001 bcd_in2=10010010 cout=1 sum=01100011
* bcd_in1=01110001 bcd_in2=10010011 cout=1 sum=01100100
* bcd_in1=01110001 bcd_in2=10010100 cout=1 sum=01100101
* bcd_in1=01110001 bcd_in2=10010101 cout=1 sum=01100110
* bcd_in1=01110001 bcd_in2=10010110 cout=1 sum=01100111
* bcd_in1=01110001 bcd_in2=10010111 cout=1 sum=01101000
* bcd_in1=01110001 bcd_in2=10011000 cout=1 sum=01101001
* bcd_in1=01110001 bcd_in2=10011001 cout=1 sum=01110000
* bcd_in1=01110010 bcd_in2=00000000 cout=0 sum=01110010
* bcd_in1=01110010 bcd_in2=00000001 cout=0 sum=01110011
* bcd_in1=01110010 bcd_in2=00000010 cout=0 sum=01110100
* bcd_in1=01110010 bcd_in2=00000011 cout=0 sum=01110101
* bcd_in1=01110010 bcd_in2=00000100 cout=0 sum=01110110
* bcd_in1=01110010 bcd_in2=00000101 cout=0 sum=01110111
* bcd_in1=01110010 bcd_in2=00000110 cout=0 sum=01111000
* bcd_in1=01110010 bcd_in2=00000111 cout=0 sum=01111001
* bcd_in1=01110010 bcd_in2=00001000 cout=0 sum=10000000
* bcd_in1=01110010 bcd_in2=00001001 cout=0 sum=10000001
* bcd_in1=01110010 bcd_in2=00010000 cout=0 sum=10000010
* bcd_in1=01110010 bcd_in2=00010001 cout=0 sum=10000011
* bcd_in1=01110010 bcd_in2=00010010 cout=0 sum=10000100
* bcd_in1=01110010 bcd_in2=00010011 cout=0 sum=10000101
* bcd_in1=01110010 bcd_in2=00010100 cout=0 sum=10000110
* bcd_in1=01110010 bcd_in2=00010101 cout=0 sum=10000111
* bcd_in1=01110010 bcd_in2=00010110 cout=0 sum=10001000
* bcd_in1=01110010 bcd_in2=00010111 cout=0 sum=10001001
* bcd_in1=01110010 bcd_in2=00011000 cout=0 sum=10010000
* bcd_in1=01110010 bcd_in2=00011001 cout=0 sum=10010001
* bcd_in1=01110010 bcd_in2=00100000 cout=0 sum=10010010
* bcd_in1=01110010 bcd_in2=00100001 cout=0 sum=10010011
* bcd_in1=01110010 bcd_in2=00100010 cout=0 sum=10010100
* bcd_in1=01110010 bcd_in2=00100011 cout=0 sum=10010101
* bcd_in1=01110010 bcd_in2=00100100 cout=0 sum=10010110
* bcd_in1=01110010 bcd_in2=00100101 cout=0 sum=10010111
* bcd_in1=01110010 bcd_in2=00100110 cout=0 sum=10011000
* bcd_in1=01110010 bcd_in2=00100111 cout=0 sum=10011001
* bcd_in1=01110010 bcd_in2=00101000 cout=1 sum=00000000
* bcd_in1=01110010 bcd_in2=00101001 cout=1 sum=00000001
* bcd_in1=01110010 bcd_in2=00110000 cout=1 sum=00000010
* bcd_in1=01110010 bcd_in2=00110001 cout=1 sum=00000011
* bcd_in1=01110010 bcd_in2=00110010 cout=1 sum=00000100
* bcd_in1=01110010 bcd_in2=00110011 cout=1 sum=00000101
* bcd_in1=01110010 bcd_in2=00110100 cout=1 sum=00000110
* bcd_in1=01110010 bcd_in2=00110101 cout=1 sum=00000111
* bcd_in1=01110010 bcd_in2=00110110 cout=1 sum=00001000
* bcd_in1=01110010 bcd_in2=00110111 cout=1 sum=00001001
* bcd_in1=01110010 bcd_in2=00111000 cout=1 sum=00010000
* bcd_in1=01110010 bcd_in2=00111001 cout=1 sum=00010001
* bcd_in1=01110010 bcd_in2=01000000 cout=1 sum=00010010
* bcd_in1=01110010 bcd_in2=01000001 cout=1 sum=00010011
* bcd_in1=01110010 bcd_in2=01000010 cout=1 sum=00010100
* bcd_in1=01110010 bcd_in2=01000011 cout=1 sum=00010101
* bcd_in1=01110010 bcd_in2=01000100 cout=1 sum=00010110
* bcd_in1=01110010 bcd_in2=01000101 cout=1 sum=00010111
* bcd_in1=01110010 bcd_in2=01000110 cout=1 sum=00011000
* bcd_in1=01110010 bcd_in2=01000111 cout=1 sum=00011001
* bcd_in1=01110010 bcd_in2=01001000 cout=1 sum=00100000
* bcd_in1=01110010 bcd_in2=01001001 cout=1 sum=00100001
* bcd_in1=01110010 bcd_in2=01010000 cout=1 sum=00100010
* bcd_in1=01110010 bcd_in2=01010001 cout=1 sum=00100011
* bcd_in1=01110010 bcd_in2=01010010 cout=1 sum=00100100
* bcd_in1=01110010 bcd_in2=01010011 cout=1 sum=00100101
* bcd_in1=01110010 bcd_in2=01010100 cout=1 sum=00100110
* bcd_in1=01110010 bcd_in2=01010101 cout=1 sum=00100111
* bcd_in1=01110010 bcd_in2=01010110 cout=1 sum=00101000
* bcd_in1=01110010 bcd_in2=01010111 cout=1 sum=00101001
* bcd_in1=01110010 bcd_in2=01011000 cout=1 sum=00110000
* bcd_in1=01110010 bcd_in2=01011001 cout=1 sum=00110001
* bcd_in1=01110010 bcd_in2=01100000 cout=1 sum=00110010
* bcd_in1=01110010 bcd_in2=01100001 cout=1 sum=00110011
* bcd_in1=01110010 bcd_in2=01100010 cout=1 sum=00110100
* bcd_in1=01110010 bcd_in2=01100011 cout=1 sum=00110101
* bcd_in1=01110010 bcd_in2=01100100 cout=1 sum=00110110
* bcd_in1=01110010 bcd_in2=01100101 cout=1 sum=00110111
* bcd_in1=01110010 bcd_in2=01100110 cout=1 sum=00111000
* bcd_in1=01110010 bcd_in2=01100111 cout=1 sum=00111001
* bcd_in1=01110010 bcd_in2=01101000 cout=1 sum=01000000
* bcd_in1=01110010 bcd_in2=01101001 cout=1 sum=01000001
* bcd_in1=01110010 bcd_in2=01110000 cout=1 sum=01000010
* bcd_in1=01110010 bcd_in2=01110001 cout=1 sum=01000011
* bcd_in1=01110010 bcd_in2=01110010 cout=1 sum=01000100
* bcd_in1=01110010 bcd_in2=01110011 cout=1 sum=01000101
* bcd_in1=01110010 bcd_in2=01110100 cout=1 sum=01000110
* bcd_in1=01110010 bcd_in2=01110101 cout=1 sum=01000111
* bcd_in1=01110010 bcd_in2=01110110 cout=1 sum=01001000
* bcd_in1=01110010 bcd_in2=01110111 cout=1 sum=01001001
* bcd_in1=01110010 bcd_in2=01111000 cout=1 sum=01010000
* bcd_in1=01110010 bcd_in2=01111001 cout=1 sum=01010001
* bcd_in1=01110010 bcd_in2=10000000 cout=1 sum=01010010
* bcd_in1=01110010 bcd_in2=10000001 cout=1 sum=01010011
* bcd_in1=01110010 bcd_in2=10000010 cout=1 sum=01010100
* bcd_in1=01110010 bcd_in2=10000011 cout=1 sum=01010101
* bcd_in1=01110010 bcd_in2=10000100 cout=1 sum=01010110
* bcd_in1=01110010 bcd_in2=10000101 cout=1 sum=01010111
* bcd_in1=01110010 bcd_in2=10000110 cout=1 sum=01011000
* bcd_in1=01110010 bcd_in2=10000111 cout=1 sum=01011001
* bcd_in1=01110010 bcd_in2=10001000 cout=1 sum=01100000
* bcd_in1=01110010 bcd_in2=10001001 cout=1 sum=01100001
* bcd_in1=01110010 bcd_in2=10010000 cout=1 sum=01100010
* bcd_in1=01110010 bcd_in2=10010001 cout=1 sum=01100011
* bcd_in1=01110010 bcd_in2=10010010 cout=1 sum=01100100
* bcd_in1=01110010 bcd_in2=10010011 cout=1 sum=01100101
* bcd_in1=01110010 bcd_in2=10010100 cout=1 sum=01100110
* bcd_in1=01110010 bcd_in2=10010101 cout=1 sum=01100111
* bcd_in1=01110010 bcd_in2=10010110 cout=1 sum=01101000
* bcd_in1=01110010 bcd_in2=10010111 cout=1 sum=01101001
* bcd_in1=01110010 bcd_in2=10011000 cout=1 sum=01110000
* bcd_in1=01110010 bcd_in2=10011001 cout=1 sum=01110001
* bcd_in1=01110011 bcd_in2=00000000 cout=0 sum=01110011
* bcd_in1=01110011 bcd_in2=00000001 cout=0 sum=01110100
* bcd_in1=01110011 bcd_in2=00000010 cout=0 sum=01110101
* bcd_in1=01110011 bcd_in2=00000011 cout=0 sum=01110110
* bcd_in1=01110011 bcd_in2=00000100 cout=0 sum=01110111
* bcd_in1=01110011 bcd_in2=00000101 cout=0 sum=01111000
* bcd_in1=01110011 bcd_in2=00000110 cout=0 sum=01111001
* bcd_in1=01110011 bcd_in2=00000111 cout=0 sum=10000000
* bcd_in1=01110011 bcd_in2=00001000 cout=0 sum=10000001
* bcd_in1=01110011 bcd_in2=00001001 cout=0 sum=10000010
* bcd_in1=01110011 bcd_in2=00010000 cout=0 sum=10000011
* bcd_in1=01110011 bcd_in2=00010001 cout=0 sum=10000100
* bcd_in1=01110011 bcd_in2=00010010 cout=0 sum=10000101
* bcd_in1=01110011 bcd_in2=00010011 cout=0 sum=10000110
* bcd_in1=01110011 bcd_in2=00010100 cout=0 sum=10000111
* bcd_in1=01110011 bcd_in2=00010101 cout=0 sum=10001000
* bcd_in1=01110011 bcd_in2=00010110 cout=0 sum=10001001
* bcd_in1=01110011 bcd_in2=00010111 cout=0 sum=10010000
* bcd_in1=01110011 bcd_in2=00011000 cout=0 sum=10010001
* bcd_in1=01110011 bcd_in2=00011001 cout=0 sum=10010010
* bcd_in1=01110011 bcd_in2=00100000 cout=0 sum=10010011
* bcd_in1=01110011 bcd_in2=00100001 cout=0 sum=10010100
* bcd_in1=01110011 bcd_in2=00100010 cout=0 sum=10010101
* bcd_in1=01110011 bcd_in2=00100011 cout=0 sum=10010110
* bcd_in1=01110011 bcd_in2=00100100 cout=0 sum=10010111
* bcd_in1=01110011 bcd_in2=00100101 cout=0 sum=10011000
* bcd_in1=01110011 bcd_in2=00100110 cout=0 sum=10011001
* bcd_in1=01110011 bcd_in2=00100111 cout=1 sum=00000000
* bcd_in1=01110011 bcd_in2=00101000 cout=1 sum=00000001
* bcd_in1=01110011 bcd_in2=00101001 cout=1 sum=00000010
* bcd_in1=01110011 bcd_in2=00110000 cout=1 sum=00000011
* bcd_in1=01110011 bcd_in2=00110001 cout=1 sum=00000100
* bcd_in1=01110011 bcd_in2=00110010 cout=1 sum=00000101
* bcd_in1=01110011 bcd_in2=00110011 cout=1 sum=00000110
* bcd_in1=01110011 bcd_in2=00110100 cout=1 sum=00000111
* bcd_in1=01110011 bcd_in2=00110101 cout=1 sum=00001000
* bcd_in1=01110011 bcd_in2=00110110 cout=1 sum=00001001
* bcd_in1=01110011 bcd_in2=00110111 cout=1 sum=00010000
* bcd_in1=01110011 bcd_in2=00111000 cout=1 sum=00010001
* bcd_in1=01110011 bcd_in2=00111001 cout=1 sum=00010010
* bcd_in1=01110011 bcd_in2=01000000 cout=1 sum=00010011
* bcd_in1=01110011 bcd_in2=01000001 cout=1 sum=00010100
* bcd_in1=01110011 bcd_in2=01000010 cout=1 sum=00010101
* bcd_in1=01110011 bcd_in2=01000011 cout=1 sum=00010110
* bcd_in1=01110011 bcd_in2=01000100 cout=1 sum=00010111
* bcd_in1=01110011 bcd_in2=01000101 cout=1 sum=00011000
* bcd_in1=01110011 bcd_in2=01000110 cout=1 sum=00011001
* bcd_in1=01110011 bcd_in2=01000111 cout=1 sum=00100000
* bcd_in1=01110011 bcd_in2=01001000 cout=1 sum=00100001
* bcd_in1=01110011 bcd_in2=01001001 cout=1 sum=00100010
* bcd_in1=01110011 bcd_in2=01010000 cout=1 sum=00100011
* bcd_in1=01110011 bcd_in2=01010001 cout=1 sum=00100100
* bcd_in1=01110011 bcd_in2=01010010 cout=1 sum=00100101
* bcd_in1=01110011 bcd_in2=01010011 cout=1 sum=00100110
* bcd_in1=01110011 bcd_in2=01010100 cout=1 sum=00100111
* bcd_in1=01110011 bcd_in2=01010101 cout=1 sum=00101000
* bcd_in1=01110011 bcd_in2=01010110 cout=1 sum=00101001
* bcd_in1=01110011 bcd_in2=01010111 cout=1 sum=00110000
* bcd_in1=01110011 bcd_in2=01011000 cout=1 sum=00110001
* bcd_in1=01110011 bcd_in2=01011001 cout=1 sum=00110010
* bcd_in1=01110011 bcd_in2=01100000 cout=1 sum=00110011
* bcd_in1=01110011 bcd_in2=01100001 cout=1 sum=00110100
* bcd_in1=01110011 bcd_in2=01100010 cout=1 sum=00110101
* bcd_in1=01110011 bcd_in2=01100011 cout=1 sum=00110110
* bcd_in1=01110011 bcd_in2=01100100 cout=1 sum=00110111
* bcd_in1=01110011 bcd_in2=01100101 cout=1 sum=00111000
* bcd_in1=01110011 bcd_in2=01100110 cout=1 sum=00111001
* bcd_in1=01110011 bcd_in2=01100111 cout=1 sum=01000000
* bcd_in1=01110011 bcd_in2=01101000 cout=1 sum=01000001
* bcd_in1=01110011 bcd_in2=01101001 cout=1 sum=01000010
* bcd_in1=01110011 bcd_in2=01110000 cout=1 sum=01000011
* bcd_in1=01110011 bcd_in2=01110001 cout=1 sum=01000100
* bcd_in1=01110011 bcd_in2=01110010 cout=1 sum=01000101
* bcd_in1=01110011 bcd_in2=01110011 cout=1 sum=01000110
* bcd_in1=01110011 bcd_in2=01110100 cout=1 sum=01000111
* bcd_in1=01110011 bcd_in2=01110101 cout=1 sum=01001000
* bcd_in1=01110011 bcd_in2=01110110 cout=1 sum=01001001
* bcd_in1=01110011 bcd_in2=01110111 cout=1 sum=01010000
* bcd_in1=01110011 bcd_in2=01111000 cout=1 sum=01010001
* bcd_in1=01110011 bcd_in2=01111001 cout=1 sum=01010010
* bcd_in1=01110011 bcd_in2=10000000 cout=1 sum=01010011
* bcd_in1=01110011 bcd_in2=10000001 cout=1 sum=01010100
* bcd_in1=01110011 bcd_in2=10000010 cout=1 sum=01010101
* bcd_in1=01110011 bcd_in2=10000011 cout=1 sum=01010110
* bcd_in1=01110011 bcd_in2=10000100 cout=1 sum=01010111
* bcd_in1=01110011 bcd_in2=10000101 cout=1 sum=01011000
* bcd_in1=01110011 bcd_in2=10000110 cout=1 sum=01011001
* bcd_in1=01110011 bcd_in2=10000111 cout=1 sum=01100000
* bcd_in1=01110011 bcd_in2=10001000 cout=1 sum=01100001
* bcd_in1=01110011 bcd_in2=10001001 cout=1 sum=01100010
* bcd_in1=01110011 bcd_in2=10010000 cout=1 sum=01100011
* bcd_in1=01110011 bcd_in2=10010001 cout=1 sum=01100100
* bcd_in1=01110011 bcd_in2=10010010 cout=1 sum=01100101
* bcd_in1=01110011 bcd_in2=10010011 cout=1 sum=01100110
* bcd_in1=01110011 bcd_in2=10010100 cout=1 sum=01100111
* bcd_in1=01110011 bcd_in2=10010101 cout=1 sum=01101000
* bcd_in1=01110011 bcd_in2=10010110 cout=1 sum=01101001
* bcd_in1=01110011 bcd_in2=10010111 cout=1 sum=01110000
* bcd_in1=01110011 bcd_in2=10011000 cout=1 sum=01110001
* bcd_in1=01110011 bcd_in2=10011001 cout=1 sum=01110010
* bcd_in1=01110100 bcd_in2=00000000 cout=0 sum=01110100
* bcd_in1=01110100 bcd_in2=00000001 cout=0 sum=01110101
* bcd_in1=01110100 bcd_in2=00000010 cout=0 sum=01110110
* bcd_in1=01110100 bcd_in2=00000011 cout=0 sum=01110111
* bcd_in1=01110100 bcd_in2=00000100 cout=0 sum=01111000
* bcd_in1=01110100 bcd_in2=00000101 cout=0 sum=01111001
* bcd_in1=01110100 bcd_in2=00000110 cout=0 sum=10000000
* bcd_in1=01110100 bcd_in2=00000111 cout=0 sum=10000001
* bcd_in1=01110100 bcd_in2=00001000 cout=0 sum=10000010
* bcd_in1=01110100 bcd_in2=00001001 cout=0 sum=10000011
* bcd_in1=01110100 bcd_in2=00010000 cout=0 sum=10000100
* bcd_in1=01110100 bcd_in2=00010001 cout=0 sum=10000101
* bcd_in1=01110100 bcd_in2=00010010 cout=0 sum=10000110
* bcd_in1=01110100 bcd_in2=00010011 cout=0 sum=10000111
* bcd_in1=01110100 bcd_in2=00010100 cout=0 sum=10001000
* bcd_in1=01110100 bcd_in2=00010101 cout=0 sum=10001001
* bcd_in1=01110100 bcd_in2=00010110 cout=0 sum=10010000
* bcd_in1=01110100 bcd_in2=00010111 cout=0 sum=10010001
* bcd_in1=01110100 bcd_in2=00011000 cout=0 sum=10010010
* bcd_in1=01110100 bcd_in2=00011001 cout=0 sum=10010011
* bcd_in1=01110100 bcd_in2=00100000 cout=0 sum=10010100
* bcd_in1=01110100 bcd_in2=00100001 cout=0 sum=10010101
* bcd_in1=01110100 bcd_in2=00100010 cout=0 sum=10010110
* bcd_in1=01110100 bcd_in2=00100011 cout=0 sum=10010111
* bcd_in1=01110100 bcd_in2=00100100 cout=0 sum=10011000
* bcd_in1=01110100 bcd_in2=00100101 cout=0 sum=10011001
* bcd_in1=01110100 bcd_in2=00100110 cout=1 sum=00000000
* bcd_in1=01110100 bcd_in2=00100111 cout=1 sum=00000001
* bcd_in1=01110100 bcd_in2=00101000 cout=1 sum=00000010
* bcd_in1=01110100 bcd_in2=00101001 cout=1 sum=00000011
* bcd_in1=01110100 bcd_in2=00110000 cout=1 sum=00000100
* bcd_in1=01110100 bcd_in2=00110001 cout=1 sum=00000101
* bcd_in1=01110100 bcd_in2=00110010 cout=1 sum=00000110
* bcd_in1=01110100 bcd_in2=00110011 cout=1 sum=00000111
* bcd_in1=01110100 bcd_in2=00110100 cout=1 sum=00001000
* bcd_in1=01110100 bcd_in2=00110101 cout=1 sum=00001001
* bcd_in1=01110100 bcd_in2=00110110 cout=1 sum=00010000
* bcd_in1=01110100 bcd_in2=00110111 cout=1 sum=00010001
* bcd_in1=01110100 bcd_in2=00111000 cout=1 sum=00010010
* bcd_in1=01110100 bcd_in2=00111001 cout=1 sum=00010011
* bcd_in1=01110100 bcd_in2=01000000 cout=1 sum=00010100
* bcd_in1=01110100 bcd_in2=01000001 cout=1 sum=00010101
* bcd_in1=01110100 bcd_in2=01000010 cout=1 sum=00010110
* bcd_in1=01110100 bcd_in2=01000011 cout=1 sum=00010111
* bcd_in1=01110100 bcd_in2=01000100 cout=1 sum=00011000
* bcd_in1=01110100 bcd_in2=01000101 cout=1 sum=00011001
* bcd_in1=01110100 bcd_in2=01000110 cout=1 sum=00100000
* bcd_in1=01110100 bcd_in2=01000111 cout=1 sum=00100001
* bcd_in1=01110100 bcd_in2=01001000 cout=1 sum=00100010
* bcd_in1=01110100 bcd_in2=01001001 cout=1 sum=00100011
* bcd_in1=01110100 bcd_in2=01010000 cout=1 sum=00100100
* bcd_in1=01110100 bcd_in2=01010001 cout=1 sum=00100101
* bcd_in1=01110100 bcd_in2=01010010 cout=1 sum=00100110
* bcd_in1=01110100 bcd_in2=01010011 cout=1 sum=00100111
* bcd_in1=01110100 bcd_in2=01010100 cout=1 sum=00101000
* bcd_in1=01110100 bcd_in2=01010101 cout=1 sum=00101001
* bcd_in1=01110100 bcd_in2=01010110 cout=1 sum=00110000
* bcd_in1=01110100 bcd_in2=01010111 cout=1 sum=00110001
* bcd_in1=01110100 bcd_in2=01011000 cout=1 sum=00110010
* bcd_in1=01110100 bcd_in2=01011001 cout=1 sum=00110011
* bcd_in1=01110100 bcd_in2=01100000 cout=1 sum=00110100
* bcd_in1=01110100 bcd_in2=01100001 cout=1 sum=00110101
* bcd_in1=01110100 bcd_in2=01100010 cout=1 sum=00110110
* bcd_in1=01110100 bcd_in2=01100011 cout=1 sum=00110111
* bcd_in1=01110100 bcd_in2=01100100 cout=1 sum=00111000
* bcd_in1=01110100 bcd_in2=01100101 cout=1 sum=00111001
* bcd_in1=01110100 bcd_in2=01100110 cout=1 sum=01000000
* bcd_in1=01110100 bcd_in2=01100111 cout=1 sum=01000001
* bcd_in1=01110100 bcd_in2=01101000 cout=1 sum=01000010
* bcd_in1=01110100 bcd_in2=01101001 cout=1 sum=01000011
* bcd_in1=01110100 bcd_in2=01110000 cout=1 sum=01000100
* bcd_in1=01110100 bcd_in2=01110001 cout=1 sum=01000101
* bcd_in1=01110100 bcd_in2=01110010 cout=1 sum=01000110
* bcd_in1=01110100 bcd_in2=01110011 cout=1 sum=01000111
* bcd_in1=01110100 bcd_in2=01110100 cout=1 sum=01001000
* bcd_in1=01110100 bcd_in2=01110101 cout=1 sum=01001001
* bcd_in1=01110100 bcd_in2=01110110 cout=1 sum=01010000
* bcd_in1=01110100 bcd_in2=01110111 cout=1 sum=01010001
* bcd_in1=01110100 bcd_in2=01111000 cout=1 sum=01010010
* bcd_in1=01110100 bcd_in2=01111001 cout=1 sum=01010011
* bcd_in1=01110100 bcd_in2=10000000 cout=1 sum=01010100
* bcd_in1=01110100 bcd_in2=10000001 cout=1 sum=01010101
* bcd_in1=01110100 bcd_in2=10000010 cout=1 sum=01010110
* bcd_in1=01110100 bcd_in2=10000011 cout=1 sum=01010111
* bcd_in1=01110100 bcd_in2=10000100 cout=1 sum=01011000
* bcd_in1=01110100 bcd_in2=10000101 cout=1 sum=01011001
* bcd_in1=01110100 bcd_in2=10000110 cout=1 sum=01100000
* bcd_in1=01110100 bcd_in2=10000111 cout=1 sum=01100001
* bcd_in1=01110100 bcd_in2=10001000 cout=1 sum=01100010
* bcd_in1=01110100 bcd_in2=10001001 cout=1 sum=01100011
* bcd_in1=01110100 bcd_in2=10010000 cout=1 sum=01100100
* bcd_in1=01110100 bcd_in2=10010001 cout=1 sum=01100101
* bcd_in1=01110100 bcd_in2=10010010 cout=1 sum=01100110
* bcd_in1=01110100 bcd_in2=10010011 cout=1 sum=01100111
* bcd_in1=01110100 bcd_in2=10010100 cout=1 sum=01101000
* bcd_in1=01110100 bcd_in2=10010101 cout=1 sum=01101001
* bcd_in1=01110100 bcd_in2=10010110 cout=1 sum=01110000
* bcd_in1=01110100 bcd_in2=10010111 cout=1 sum=01110001
* bcd_in1=01110100 bcd_in2=10011000 cout=1 sum=01110010
* bcd_in1=01110100 bcd_in2=10011001 cout=1 sum=01110011
* bcd_in1=01110101 bcd_in2=00000000 cout=0 sum=01110101
* bcd_in1=01110101 bcd_in2=00000001 cout=0 sum=01110110
* bcd_in1=01110101 bcd_in2=00000010 cout=0 sum=01110111
* bcd_in1=01110101 bcd_in2=00000011 cout=0 sum=01111000
* bcd_in1=01110101 bcd_in2=00000100 cout=0 sum=01111001
* bcd_in1=01110101 bcd_in2=00000101 cout=0 sum=10000000
* bcd_in1=01110101 bcd_in2=00000110 cout=0 sum=10000001
* bcd_in1=01110101 bcd_in2=00000111 cout=0 sum=10000010
* bcd_in1=01110101 bcd_in2=00001000 cout=0 sum=10000011
* bcd_in1=01110101 bcd_in2=00001001 cout=0 sum=10000100
* bcd_in1=01110101 bcd_in2=00010000 cout=0 sum=10000101
* bcd_in1=01110101 bcd_in2=00010001 cout=0 sum=10000110
* bcd_in1=01110101 bcd_in2=00010010 cout=0 sum=10000111
* bcd_in1=01110101 bcd_in2=00010011 cout=0 sum=10001000
* bcd_in1=01110101 bcd_in2=00010100 cout=0 sum=10001001
* bcd_in1=01110101 bcd_in2=00010101 cout=0 sum=10010000
* bcd_in1=01110101 bcd_in2=00010110 cout=0 sum=10010001
* bcd_in1=01110101 bcd_in2=00010111 cout=0 sum=10010010
* bcd_in1=01110101 bcd_in2=00011000 cout=0 sum=10010011
* bcd_in1=01110101 bcd_in2=00011001 cout=0 sum=10010100
* bcd_in1=01110101 bcd_in2=00100000 cout=0 sum=10010101
* bcd_in1=01110101 bcd_in2=00100001 cout=0 sum=10010110
* bcd_in1=01110101 bcd_in2=00100010 cout=0 sum=10010111
* bcd_in1=01110101 bcd_in2=00100011 cout=0 sum=10011000
* bcd_in1=01110101 bcd_in2=00100100 cout=0 sum=10011001
* bcd_in1=01110101 bcd_in2=00100101 cout=1 sum=00000000
* bcd_in1=01110101 bcd_in2=00100110 cout=1 sum=00000001
* bcd_in1=01110101 bcd_in2=00100111 cout=1 sum=00000010
* bcd_in1=01110101 bcd_in2=00101000 cout=1 sum=00000011
* bcd_in1=01110101 bcd_in2=00101001 cout=1 sum=00000100
* bcd_in1=01110101 bcd_in2=00110000 cout=1 sum=00000101
* bcd_in1=01110101 bcd_in2=00110001 cout=1 sum=00000110
* bcd_in1=01110101 bcd_in2=00110010 cout=1 sum=00000111
* bcd_in1=01110101 bcd_in2=00110011 cout=1 sum=00001000
* bcd_in1=01110101 bcd_in2=00110100 cout=1 sum=00001001
* bcd_in1=01110101 bcd_in2=00110101 cout=1 sum=00010000
* bcd_in1=01110101 bcd_in2=00110110 cout=1 sum=00010001
* bcd_in1=01110101 bcd_in2=00110111 cout=1 sum=00010010
* bcd_in1=01110101 bcd_in2=00111000 cout=1 sum=00010011
* bcd_in1=01110101 bcd_in2=00111001 cout=1 sum=00010100
* bcd_in1=01110101 bcd_in2=01000000 cout=1 sum=00010101
* bcd_in1=01110101 bcd_in2=01000001 cout=1 sum=00010110
* bcd_in1=01110101 bcd_in2=01000010 cout=1 sum=00010111
* bcd_in1=01110101 bcd_in2=01000011 cout=1 sum=00011000
* bcd_in1=01110101 bcd_in2=01000100 cout=1 sum=00011001
* bcd_in1=01110101 bcd_in2=01000101 cout=1 sum=00100000
* bcd_in1=01110101 bcd_in2=01000110 cout=1 sum=00100001
* bcd_in1=01110101 bcd_in2=01000111 cout=1 sum=00100010
* bcd_in1=01110101 bcd_in2=01001000 cout=1 sum=00100011
* bcd_in1=01110101 bcd_in2=01001001 cout=1 sum=00100100
* bcd_in1=01110101 bcd_in2=01010000 cout=1 sum=00100101
* bcd_in1=01110101 bcd_in2=01010001 cout=1 sum=00100110
* bcd_in1=01110101 bcd_in2=01010010 cout=1 sum=00100111
* bcd_in1=01110101 bcd_in2=01010011 cout=1 sum=00101000
* bcd_in1=01110101 bcd_in2=01010100 cout=1 sum=00101001
* bcd_in1=01110101 bcd_in2=01010101 cout=1 sum=00110000
* bcd_in1=01110101 bcd_in2=01010110 cout=1 sum=00110001
* bcd_in1=01110101 bcd_in2=01010111 cout=1 sum=00110010
* bcd_in1=01110101 bcd_in2=01011000 cout=1 sum=00110011
* bcd_in1=01110101 bcd_in2=01011001 cout=1 sum=00110100
* bcd_in1=01110101 bcd_in2=01100000 cout=1 sum=00110101
* bcd_in1=01110101 bcd_in2=01100001 cout=1 sum=00110110
* bcd_in1=01110101 bcd_in2=01100010 cout=1 sum=00110111
* bcd_in1=01110101 bcd_in2=01100011 cout=1 sum=00111000
* bcd_in1=01110101 bcd_in2=01100100 cout=1 sum=00111001
* bcd_in1=01110101 bcd_in2=01100101 cout=1 sum=01000000
* bcd_in1=01110101 bcd_in2=01100110 cout=1 sum=01000001
* bcd_in1=01110101 bcd_in2=01100111 cout=1 sum=01000010
* bcd_in1=01110101 bcd_in2=01101000 cout=1 sum=01000011
* bcd_in1=01110101 bcd_in2=01101001 cout=1 sum=01000100
* bcd_in1=01110101 bcd_in2=01110000 cout=1 sum=01000101
* bcd_in1=01110101 bcd_in2=01110001 cout=1 sum=01000110
* bcd_in1=01110101 bcd_in2=01110010 cout=1 sum=01000111
* bcd_in1=01110101 bcd_in2=01110011 cout=1 sum=01001000
* bcd_in1=01110101 bcd_in2=01110100 cout=1 sum=01001001
* bcd_in1=01110101 bcd_in2=01110101 cout=1 sum=01010000
* bcd_in1=01110101 bcd_in2=01110110 cout=1 sum=01010001
* bcd_in1=01110101 bcd_in2=01110111 cout=1 sum=01010010
* bcd_in1=01110101 bcd_in2=01111000 cout=1 sum=01010011
* bcd_in1=01110101 bcd_in2=01111001 cout=1 sum=01010100
* bcd_in1=01110101 bcd_in2=10000000 cout=1 sum=01010101
* bcd_in1=01110101 bcd_in2=10000001 cout=1 sum=01010110
* bcd_in1=01110101 bcd_in2=10000010 cout=1 sum=01010111
* bcd_in1=01110101 bcd_in2=10000011 cout=1 sum=01011000
* bcd_in1=01110101 bcd_in2=10000100 cout=1 sum=01011001
* bcd_in1=01110101 bcd_in2=10000101 cout=1 sum=01100000
* bcd_in1=01110101 bcd_in2=10000110 cout=1 sum=01100001
* bcd_in1=01110101 bcd_in2=10000111 cout=1 sum=01100010
* bcd_in1=01110101 bcd_in2=10001000 cout=1 sum=01100011
* bcd_in1=01110101 bcd_in2=10001001 cout=1 sum=01100100
* bcd_in1=01110101 bcd_in2=10010000 cout=1 sum=01100101
* bcd_in1=01110101 bcd_in2=10010001 cout=1 sum=01100110
* bcd_in1=01110101 bcd_in2=10010010 cout=1 sum=01100111
* bcd_in1=01110101 bcd_in2=10010011 cout=1 sum=01101000
* bcd_in1=01110101 bcd_in2=10010100 cout=1 sum=01101001
* bcd_in1=01110101 bcd_in2=10010101 cout=1 sum=01110000
* bcd_in1=01110101 bcd_in2=10010110 cout=1 sum=01110001
* bcd_in1=01110101 bcd_in2=10010111 cout=1 sum=01110010
* bcd_in1=01110101 bcd_in2=10011000 cout=1 sum=01110011
* bcd_in1=01110101 bcd_in2=10011001 cout=1 sum=01110100
* bcd_in1=01110110 bcd_in2=00000000 cout=0 sum=01110110
* bcd_in1=01110110 bcd_in2=00000001 cout=0 sum=01110111
* bcd_in1=01110110 bcd_in2=00000010 cout=0 sum=01111000
* bcd_in1=01110110 bcd_in2=00000011 cout=0 sum=01111001
* bcd_in1=01110110 bcd_in2=00000100 cout=0 sum=10000000
* bcd_in1=01110110 bcd_in2=00000101 cout=0 sum=10000001
* bcd_in1=01110110 bcd_in2=00000110 cout=0 sum=10000010
* bcd_in1=01110110 bcd_in2=00000111 cout=0 sum=10000011
* bcd_in1=01110110 bcd_in2=00001000 cout=0 sum=10000100
* bcd_in1=01110110 bcd_in2=00001001 cout=0 sum=10000101
* bcd_in1=01110110 bcd_in2=00010000 cout=0 sum=10000110
* bcd_in1=01110110 bcd_in2=00010001 cout=0 sum=10000111
* bcd_in1=01110110 bcd_in2=00010010 cout=0 sum=10001000
* bcd_in1=01110110 bcd_in2=00010011 cout=0 sum=10001001
* bcd_in1=01110110 bcd_in2=00010100 cout=0 sum=10010000
* bcd_in1=01110110 bcd_in2=00010101 cout=0 sum=10010001
* bcd_in1=01110110 bcd_in2=00010110 cout=0 sum=10010010
* bcd_in1=01110110 bcd_in2=00010111 cout=0 sum=10010011
* bcd_in1=01110110 bcd_in2=00011000 cout=0 sum=10010100
* bcd_in1=01110110 bcd_in2=00011001 cout=0 sum=10010101
* bcd_in1=01110110 bcd_in2=00100000 cout=0 sum=10010110
* bcd_in1=01110110 bcd_in2=00100001 cout=0 sum=10010111
* bcd_in1=01110110 bcd_in2=00100010 cout=0 sum=10011000
* bcd_in1=01110110 bcd_in2=00100011 cout=0 sum=10011001
* bcd_in1=01110110 bcd_in2=00100100 cout=1 sum=00000000
* bcd_in1=01110110 bcd_in2=00100101 cout=1 sum=00000001
* bcd_in1=01110110 bcd_in2=00100110 cout=1 sum=00000010
* bcd_in1=01110110 bcd_in2=00100111 cout=1 sum=00000011
* bcd_in1=01110110 bcd_in2=00101000 cout=1 sum=00000100
* bcd_in1=01110110 bcd_in2=00101001 cout=1 sum=00000101
* bcd_in1=01110110 bcd_in2=00110000 cout=1 sum=00000110
* bcd_in1=01110110 bcd_in2=00110001 cout=1 sum=00000111
* bcd_in1=01110110 bcd_in2=00110010 cout=1 sum=00001000
* bcd_in1=01110110 bcd_in2=00110011 cout=1 sum=00001001
* bcd_in1=01110110 bcd_in2=00110100 cout=1 sum=00010000
* bcd_in1=01110110 bcd_in2=00110101 cout=1 sum=00010001
* bcd_in1=01110110 bcd_in2=00110110 cout=1 sum=00010010
* bcd_in1=01110110 bcd_in2=00110111 cout=1 sum=00010011
* bcd_in1=01110110 bcd_in2=00111000 cout=1 sum=00010100
* bcd_in1=01110110 bcd_in2=00111001 cout=1 sum=00010101
* bcd_in1=01110110 bcd_in2=01000000 cout=1 sum=00010110
* bcd_in1=01110110 bcd_in2=01000001 cout=1 sum=00010111
* bcd_in1=01110110 bcd_in2=01000010 cout=1 sum=00011000
* bcd_in1=01110110 bcd_in2=01000011 cout=1 sum=00011001
* bcd_in1=01110110 bcd_in2=01000100 cout=1 sum=00100000
* bcd_in1=01110110 bcd_in2=01000101 cout=1 sum=00100001
* bcd_in1=01110110 bcd_in2=01000110 cout=1 sum=00100010
* bcd_in1=01110110 bcd_in2=01000111 cout=1 sum=00100011
* bcd_in1=01110110 bcd_in2=01001000 cout=1 sum=00100100
* bcd_in1=01110110 bcd_in2=01001001 cout=1 sum=00100101
* bcd_in1=01110110 bcd_in2=01010000 cout=1 sum=00100110
* bcd_in1=01110110 bcd_in2=01010001 cout=1 sum=00100111
* bcd_in1=01110110 bcd_in2=01010010 cout=1 sum=00101000
* bcd_in1=01110110 bcd_in2=01010011 cout=1 sum=00101001
* bcd_in1=01110110 bcd_in2=01010100 cout=1 sum=00110000
* bcd_in1=01110110 bcd_in2=01010101 cout=1 sum=00110001
* bcd_in1=01110110 bcd_in2=01010110 cout=1 sum=00110010
* bcd_in1=01110110 bcd_in2=01010111 cout=1 sum=00110011
* bcd_in1=01110110 bcd_in2=01011000 cout=1 sum=00110100
* bcd_in1=01110110 bcd_in2=01011001 cout=1 sum=00110101
* bcd_in1=01110110 bcd_in2=01100000 cout=1 sum=00110110
* bcd_in1=01110110 bcd_in2=01100001 cout=1 sum=00110111
* bcd_in1=01110110 bcd_in2=01100010 cout=1 sum=00111000
* bcd_in1=01110110 bcd_in2=01100011 cout=1 sum=00111001
* bcd_in1=01110110 bcd_in2=01100100 cout=1 sum=01000000
* bcd_in1=01110110 bcd_in2=01100101 cout=1 sum=01000001
* bcd_in1=01110110 bcd_in2=01100110 cout=1 sum=01000010
* bcd_in1=01110110 bcd_in2=01100111 cout=1 sum=01000011
* bcd_in1=01110110 bcd_in2=01101000 cout=1 sum=01000100
* bcd_in1=01110110 bcd_in2=01101001 cout=1 sum=01000101
* bcd_in1=01110110 bcd_in2=01110000 cout=1 sum=01000110
* bcd_in1=01110110 bcd_in2=01110001 cout=1 sum=01000111
* bcd_in1=01110110 bcd_in2=01110010 cout=1 sum=01001000
* bcd_in1=01110110 bcd_in2=01110011 cout=1 sum=01001001
* bcd_in1=01110110 bcd_in2=01110100 cout=1 sum=01010000
* bcd_in1=01110110 bcd_in2=01110101 cout=1 sum=01010001
* bcd_in1=01110110 bcd_in2=01110110 cout=1 sum=01010010
* bcd_in1=01110110 bcd_in2=01110111 cout=1 sum=01010011
* bcd_in1=01110110 bcd_in2=01111000 cout=1 sum=01010100
* bcd_in1=01110110 bcd_in2=01111001 cout=1 sum=01010101
* bcd_in1=01110110 bcd_in2=10000000 cout=1 sum=01010110
* bcd_in1=01110110 bcd_in2=10000001 cout=1 sum=01010111
* bcd_in1=01110110 bcd_in2=10000010 cout=1 sum=01011000
* bcd_in1=01110110 bcd_in2=10000011 cout=1 sum=01011001
* bcd_in1=01110110 bcd_in2=10000100 cout=1 sum=01100000
* bcd_in1=01110110 bcd_in2=10000101 cout=1 sum=01100001
* bcd_in1=01110110 bcd_in2=10000110 cout=1 sum=01100010
* bcd_in1=01110110 bcd_in2=10000111 cout=1 sum=01100011
* bcd_in1=01110110 bcd_in2=10001000 cout=1 sum=01100100
* bcd_in1=01110110 bcd_in2=10001001 cout=1 sum=01100101
* bcd_in1=01110110 bcd_in2=10010000 cout=1 sum=01100110
* bcd_in1=01110110 bcd_in2=10010001 cout=1 sum=01100111
* bcd_in1=01110110 bcd_in2=10010010 cout=1 sum=01101000
* bcd_in1=01110110 bcd_in2=10010011 cout=1 sum=01101001
* bcd_in1=01110110 bcd_in2=10010100 cout=1 sum=01110000
* bcd_in1=01110110 bcd_in2=10010101 cout=1 sum=01110001
* bcd_in1=01110110 bcd_in2=10010110 cout=1 sum=01110010
* bcd_in1=01110110 bcd_in2=10010111 cout=1 sum=01110011
* bcd_in1=01110110 bcd_in2=10011000 cout=1 sum=01110100
* bcd_in1=01110110 bcd_in2=10011001 cout=1 sum=01110101
* bcd_in1=01110111 bcd_in2=00000000 cout=0 sum=01110111
* bcd_in1=01110111 bcd_in2=00000001 cout=0 sum=01111000
* bcd_in1=01110111 bcd_in2=00000010 cout=0 sum=01111001
* bcd_in1=01110111 bcd_in2=00000011 cout=0 sum=10000000
* bcd_in1=01110111 bcd_in2=00000100 cout=0 sum=10000001
* bcd_in1=01110111 bcd_in2=00000101 cout=0 sum=10000010
* bcd_in1=01110111 bcd_in2=00000110 cout=0 sum=10000011
* bcd_in1=01110111 bcd_in2=00000111 cout=0 sum=10000100
* bcd_in1=01110111 bcd_in2=00001000 cout=0 sum=10000101
* bcd_in1=01110111 bcd_in2=00001001 cout=0 sum=10000110
* bcd_in1=01110111 bcd_in2=00010000 cout=0 sum=10000111
* bcd_in1=01110111 bcd_in2=00010001 cout=0 sum=10001000
* bcd_in1=01110111 bcd_in2=00010010 cout=0 sum=10001001
* bcd_in1=01110111 bcd_in2=00010011 cout=0 sum=10010000
* bcd_in1=01110111 bcd_in2=00010100 cout=0 sum=10010001
* bcd_in1=01110111 bcd_in2=00010101 cout=0 sum=10010010
* bcd_in1=01110111 bcd_in2=00010110 cout=0 sum=10010011
* bcd_in1=01110111 bcd_in2=00010111 cout=0 sum=10010100
* bcd_in1=01110111 bcd_in2=00011000 cout=0 sum=10010101
* bcd_in1=01110111 bcd_in2=00011001 cout=0 sum=10010110
* bcd_in1=01110111 bcd_in2=00100000 cout=0 sum=10010111
* bcd_in1=01110111 bcd_in2=00100001 cout=0 sum=10011000
* bcd_in1=01110111 bcd_in2=00100010 cout=0 sum=10011001
* bcd_in1=01110111 bcd_in2=00100011 cout=1 sum=00000000
* bcd_in1=01110111 bcd_in2=00100100 cout=1 sum=00000001
* bcd_in1=01110111 bcd_in2=00100101 cout=1 sum=00000010
* bcd_in1=01110111 bcd_in2=00100110 cout=1 sum=00000011
* bcd_in1=01110111 bcd_in2=00100111 cout=1 sum=00000100
* bcd_in1=01110111 bcd_in2=00101000 cout=1 sum=00000101
* bcd_in1=01110111 bcd_in2=00101001 cout=1 sum=00000110
* bcd_in1=01110111 bcd_in2=00110000 cout=1 sum=00000111
* bcd_in1=01110111 bcd_in2=00110001 cout=1 sum=00001000
* bcd_in1=01110111 bcd_in2=00110010 cout=1 sum=00001001
* bcd_in1=01110111 bcd_in2=00110011 cout=1 sum=00010000
* bcd_in1=01110111 bcd_in2=00110100 cout=1 sum=00010001
* bcd_in1=01110111 bcd_in2=00110101 cout=1 sum=00010010
* bcd_in1=01110111 bcd_in2=00110110 cout=1 sum=00010011
* bcd_in1=01110111 bcd_in2=00110111 cout=1 sum=00010100
* bcd_in1=01110111 bcd_in2=00111000 cout=1 sum=00010101
* bcd_in1=01110111 bcd_in2=00111001 cout=1 sum=00010110
* bcd_in1=01110111 bcd_in2=01000000 cout=1 sum=00010111
* bcd_in1=01110111 bcd_in2=01000001 cout=1 sum=00011000
* bcd_in1=01110111 bcd_in2=01000010 cout=1 sum=00011001
* bcd_in1=01110111 bcd_in2=01000011 cout=1 sum=00100000
* bcd_in1=01110111 bcd_in2=01000100 cout=1 sum=00100001
* bcd_in1=01110111 bcd_in2=01000101 cout=1 sum=00100010
* bcd_in1=01110111 bcd_in2=01000110 cout=1 sum=00100011
* bcd_in1=01110111 bcd_in2=01000111 cout=1 sum=00100100
* bcd_in1=01110111 bcd_in2=01001000 cout=1 sum=00100101
* bcd_in1=01110111 bcd_in2=01001001 cout=1 sum=00100110
* bcd_in1=01110111 bcd_in2=01010000 cout=1 sum=00100111
* bcd_in1=01110111 bcd_in2=01010001 cout=1 sum=00101000
* bcd_in1=01110111 bcd_in2=01010010 cout=1 sum=00101001
* bcd_in1=01110111 bcd_in2=01010011 cout=1 sum=00110000
* bcd_in1=01110111 bcd_in2=01010100 cout=1 sum=00110001
* bcd_in1=01110111 bcd_in2=01010101 cout=1 sum=00110010
* bcd_in1=01110111 bcd_in2=01010110 cout=1 sum=00110011
* bcd_in1=01110111 bcd_in2=01010111 cout=1 sum=00110100
* bcd_in1=01110111 bcd_in2=01011000 cout=1 sum=00110101
* bcd_in1=01110111 bcd_in2=01011001 cout=1 sum=00110110
* bcd_in1=01110111 bcd_in2=01100000 cout=1 sum=00110111
* bcd_in1=01110111 bcd_in2=01100001 cout=1 sum=00111000
* bcd_in1=01110111 bcd_in2=01100010 cout=1 sum=00111001
* bcd_in1=01110111 bcd_in2=01100011 cout=1 sum=01000000
* bcd_in1=01110111 bcd_in2=01100100 cout=1 sum=01000001
* bcd_in1=01110111 bcd_in2=01100101 cout=1 sum=01000010
* bcd_in1=01110111 bcd_in2=01100110 cout=1 sum=01000011
* bcd_in1=01110111 bcd_in2=01100111 cout=1 sum=01000100
* bcd_in1=01110111 bcd_in2=01101000 cout=1 sum=01000101
* bcd_in1=01110111 bcd_in2=01101001 cout=1 sum=01000110
* bcd_in1=01110111 bcd_in2=01110000 cout=1 sum=01000111
* bcd_in1=01110111 bcd_in2=01110001 cout=1 sum=01001000
* bcd_in1=01110111 bcd_in2=01110010 cout=1 sum=01001001
* bcd_in1=01110111 bcd_in2=01110011 cout=1 sum=01010000
* bcd_in1=01110111 bcd_in2=01110100 cout=1 sum=01010001
* bcd_in1=01110111 bcd_in2=01110101 cout=1 sum=01010010
* bcd_in1=01110111 bcd_in2=01110110 cout=1 sum=01010011
* bcd_in1=01110111 bcd_in2=01110111 cout=1 sum=01010100
* bcd_in1=01110111 bcd_in2=01111000 cout=1 sum=01010101
* bcd_in1=01110111 bcd_in2=01111001 cout=1 sum=01010110
* bcd_in1=01110111 bcd_in2=10000000 cout=1 sum=01010111
* bcd_in1=01110111 bcd_in2=10000001 cout=1 sum=01011000
* bcd_in1=01110111 bcd_in2=10000010 cout=1 sum=01011001
* bcd_in1=01110111 bcd_in2=10000011 cout=1 sum=01100000
* bcd_in1=01110111 bcd_in2=10000100 cout=1 sum=01100001
* bcd_in1=01110111 bcd_in2=10000101 cout=1 sum=01100010
* bcd_in1=01110111 bcd_in2=10000110 cout=1 sum=01100011
* bcd_in1=01110111 bcd_in2=10000111 cout=1 sum=01100100
* bcd_in1=01110111 bcd_in2=10001000 cout=1 sum=01100101
* bcd_in1=01110111 bcd_in2=10001001 cout=1 sum=01100110
* bcd_in1=01110111 bcd_in2=10010000 cout=1 sum=01100111
* bcd_in1=01110111 bcd_in2=10010001 cout=1 sum=01101000
* bcd_in1=01110111 bcd_in2=10010010 cout=1 sum=01101001
* bcd_in1=01110111 bcd_in2=10010011 cout=1 sum=01110000
* bcd_in1=01110111 bcd_in2=10010100 cout=1 sum=01110001
* bcd_in1=01110111 bcd_in2=10010101 cout=1 sum=01110010
* bcd_in1=01110111 bcd_in2=10010110 cout=1 sum=01110011
* bcd_in1=01110111 bcd_in2=10010111 cout=1 sum=01110100
* bcd_in1=01110111 bcd_in2=10011000 cout=1 sum=01110101
* bcd_in1=01110111 bcd_in2=10011001 cout=1 sum=01110110
* bcd_in1=01111000 bcd_in2=00000000 cout=0 sum=01111000
* bcd_in1=01111000 bcd_in2=00000001 cout=0 sum=01111001
* bcd_in1=01111000 bcd_in2=00000010 cout=0 sum=10000000
* bcd_in1=01111000 bcd_in2=00000011 cout=0 sum=10000001
* bcd_in1=01111000 bcd_in2=00000100 cout=0 sum=10000010
* bcd_in1=01111000 bcd_in2=00000101 cout=0 sum=10000011
* bcd_in1=01111000 bcd_in2=00000110 cout=0 sum=10000100
* bcd_in1=01111000 bcd_in2=00000111 cout=0 sum=10000101
* bcd_in1=01111000 bcd_in2=00001000 cout=0 sum=10000110
* bcd_in1=01111000 bcd_in2=00001001 cout=0 sum=10000111
* bcd_in1=01111000 bcd_in2=00010000 cout=0 sum=10001000
* bcd_in1=01111000 bcd_in2=00010001 cout=0 sum=10001001
* bcd_in1=01111000 bcd_in2=00010010 cout=0 sum=10010000
* bcd_in1=01111000 bcd_in2=00010011 cout=0 sum=10010001
* bcd_in1=01111000 bcd_in2=00010100 cout=0 sum=10010010
* bcd_in1=01111000 bcd_in2=00010101 cout=0 sum=10010011
* bcd_in1=01111000 bcd_in2=00010110 cout=0 sum=10010100
* bcd_in1=01111000 bcd_in2=00010111 cout=0 sum=10010101
* bcd_in1=01111000 bcd_in2=00011000 cout=0 sum=10010110
* bcd_in1=01111000 bcd_in2=00011001 cout=0 sum=10010111
* bcd_in1=01111000 bcd_in2=00100000 cout=0 sum=10011000
* bcd_in1=01111000 bcd_in2=00100001 cout=0 sum=10011001
* bcd_in1=01111000 bcd_in2=00100010 cout=1 sum=00000000
* bcd_in1=01111000 bcd_in2=00100011 cout=1 sum=00000001
* bcd_in1=01111000 bcd_in2=00100100 cout=1 sum=00000010
* bcd_in1=01111000 bcd_in2=00100101 cout=1 sum=00000011
* bcd_in1=01111000 bcd_in2=00100110 cout=1 sum=00000100
* bcd_in1=01111000 bcd_in2=00100111 cout=1 sum=00000101
* bcd_in1=01111000 bcd_in2=00101000 cout=1 sum=00000110
* bcd_in1=01111000 bcd_in2=00101001 cout=1 sum=00000111
* bcd_in1=01111000 bcd_in2=00110000 cout=1 sum=00001000
* bcd_in1=01111000 bcd_in2=00110001 cout=1 sum=00001001
* bcd_in1=01111000 bcd_in2=00110010 cout=1 sum=00010000
* bcd_in1=01111000 bcd_in2=00110011 cout=1 sum=00010001
* bcd_in1=01111000 bcd_in2=00110100 cout=1 sum=00010010
* bcd_in1=01111000 bcd_in2=00110101 cout=1 sum=00010011
* bcd_in1=01111000 bcd_in2=00110110 cout=1 sum=00010100
* bcd_in1=01111000 bcd_in2=00110111 cout=1 sum=00010101
* bcd_in1=01111000 bcd_in2=00111000 cout=1 sum=00010110
* bcd_in1=01111000 bcd_in2=00111001 cout=1 sum=00010111
* bcd_in1=01111000 bcd_in2=01000000 cout=1 sum=00011000
* bcd_in1=01111000 bcd_in2=01000001 cout=1 sum=00011001
* bcd_in1=01111000 bcd_in2=01000010 cout=1 sum=00100000
* bcd_in1=01111000 bcd_in2=01000011 cout=1 sum=00100001
* bcd_in1=01111000 bcd_in2=01000100 cout=1 sum=00100010
* bcd_in1=01111000 bcd_in2=01000101 cout=1 sum=00100011
* bcd_in1=01111000 bcd_in2=01000110 cout=1 sum=00100100
* bcd_in1=01111000 bcd_in2=01000111 cout=1 sum=00100101
* bcd_in1=01111000 bcd_in2=01001000 cout=1 sum=00100110
* bcd_in1=01111000 bcd_in2=01001001 cout=1 sum=00100111
* bcd_in1=01111000 bcd_in2=01010000 cout=1 sum=00101000
* bcd_in1=01111000 bcd_in2=01010001 cout=1 sum=00101001
* bcd_in1=01111000 bcd_in2=01010010 cout=1 sum=00110000
* bcd_in1=01111000 bcd_in2=01010011 cout=1 sum=00110001
* bcd_in1=01111000 bcd_in2=01010100 cout=1 sum=00110010
* bcd_in1=01111000 bcd_in2=01010101 cout=1 sum=00110011
* bcd_in1=01111000 bcd_in2=01010110 cout=1 sum=00110100
* bcd_in1=01111000 bcd_in2=01010111 cout=1 sum=00110101
* bcd_in1=01111000 bcd_in2=01011000 cout=1 sum=00110110
* bcd_in1=01111000 bcd_in2=01011001 cout=1 sum=00110111
* bcd_in1=01111000 bcd_in2=01100000 cout=1 sum=00111000
* bcd_in1=01111000 bcd_in2=01100001 cout=1 sum=00111001
* bcd_in1=01111000 bcd_in2=01100010 cout=1 sum=01000000
* bcd_in1=01111000 bcd_in2=01100011 cout=1 sum=01000001
* bcd_in1=01111000 bcd_in2=01100100 cout=1 sum=01000010
* bcd_in1=01111000 bcd_in2=01100101 cout=1 sum=01000011
* bcd_in1=01111000 bcd_in2=01100110 cout=1 sum=01000100
* bcd_in1=01111000 bcd_in2=01100111 cout=1 sum=01000101
* bcd_in1=01111000 bcd_in2=01101000 cout=1 sum=01000110
* bcd_in1=01111000 bcd_in2=01101001 cout=1 sum=01000111
* bcd_in1=01111000 bcd_in2=01110000 cout=1 sum=01001000
* bcd_in1=01111000 bcd_in2=01110001 cout=1 sum=01001001
* bcd_in1=01111000 bcd_in2=01110010 cout=1 sum=01010000
* bcd_in1=01111000 bcd_in2=01110011 cout=1 sum=01010001
* bcd_in1=01111000 bcd_in2=01110100 cout=1 sum=01010010
* bcd_in1=01111000 bcd_in2=01110101 cout=1 sum=01010011
* bcd_in1=01111000 bcd_in2=01110110 cout=1 sum=01010100
* bcd_in1=01111000 bcd_in2=01110111 cout=1 sum=01010101
* bcd_in1=01111000 bcd_in2=01111000 cout=1 sum=01010110
* bcd_in1=01111000 bcd_in2=01111001 cout=1 sum=01010111
* bcd_in1=01111000 bcd_in2=10000000 cout=1 sum=01011000
* bcd_in1=01111000 bcd_in2=10000001 cout=1 sum=01011001
* bcd_in1=01111000 bcd_in2=10000010 cout=1 sum=01100000
* bcd_in1=01111000 bcd_in2=10000011 cout=1 sum=01100001
* bcd_in1=01111000 bcd_in2=10000100 cout=1 sum=01100010
* bcd_in1=01111000 bcd_in2=10000101 cout=1 sum=01100011
* bcd_in1=01111000 bcd_in2=10000110 cout=1 sum=01100100
* bcd_in1=01111000 bcd_in2=10000111 cout=1 sum=01100101
* bcd_in1=01111000 bcd_in2=10001000 cout=1 sum=01100110
* bcd_in1=01111000 bcd_in2=10001001 cout=1 sum=01100111
* bcd_in1=01111000 bcd_in2=10010000 cout=1 sum=01101000
* bcd_in1=01111000 bcd_in2=10010001 cout=1 sum=01101001
* bcd_in1=01111000 bcd_in2=10010010 cout=1 sum=01110000
* bcd_in1=01111000 bcd_in2=10010011 cout=1 sum=01110001
* bcd_in1=01111000 bcd_in2=10010100 cout=1 sum=01110010
* bcd_in1=01111000 bcd_in2=10010101 cout=1 sum=01110011
* bcd_in1=01111000 bcd_in2=10010110 cout=1 sum=01110100
* bcd_in1=01111000 bcd_in2=10010111 cout=1 sum=01110101
* bcd_in1=01111000 bcd_in2=10011000 cout=1 sum=01110110
* bcd_in1=01111000 bcd_in2=10011001 cout=1 sum=01110111
* bcd_in1=01111001 bcd_in2=00000000 cout=0 sum=01111001
* bcd_in1=01111001 bcd_in2=00000001 cout=0 sum=10000000
* bcd_in1=01111001 bcd_in2=00000010 cout=0 sum=10000001
* bcd_in1=01111001 bcd_in2=00000011 cout=0 sum=10000010
* bcd_in1=01111001 bcd_in2=00000100 cout=0 sum=10000011
* bcd_in1=01111001 bcd_in2=00000101 cout=0 sum=10000100
* bcd_in1=01111001 bcd_in2=00000110 cout=0 sum=10000101
* bcd_in1=01111001 bcd_in2=00000111 cout=0 sum=10000110
* bcd_in1=01111001 bcd_in2=00001000 cout=0 sum=10000111
* bcd_in1=01111001 bcd_in2=00001001 cout=0 sum=10001000
* bcd_in1=01111001 bcd_in2=00010000 cout=0 sum=10001001
* bcd_in1=01111001 bcd_in2=00010001 cout=0 sum=10010000
* bcd_in1=01111001 bcd_in2=00010010 cout=0 sum=10010001
* bcd_in1=01111001 bcd_in2=00010011 cout=0 sum=10010010
* bcd_in1=01111001 bcd_in2=00010100 cout=0 sum=10010011
* bcd_in1=01111001 bcd_in2=00010101 cout=0 sum=10010100
* bcd_in1=01111001 bcd_in2=00010110 cout=0 sum=10010101
* bcd_in1=01111001 bcd_in2=00010111 cout=0 sum=10010110
* bcd_in1=01111001 bcd_in2=00011000 cout=0 sum=10010111
* bcd_in1=01111001 bcd_in2=00011001 cout=0 sum=10011000
* bcd_in1=01111001 bcd_in2=00100000 cout=0 sum=10011001
* bcd_in1=01111001 bcd_in2=00100001 cout=1 sum=00000000
* bcd_in1=01111001 bcd_in2=00100010 cout=1 sum=00000001
* bcd_in1=01111001 bcd_in2=00100011 cout=1 sum=00000010
* bcd_in1=01111001 bcd_in2=00100100 cout=1 sum=00000011
* bcd_in1=01111001 bcd_in2=00100101 cout=1 sum=00000100
* bcd_in1=01111001 bcd_in2=00100110 cout=1 sum=00000101
* bcd_in1=01111001 bcd_in2=00100111 cout=1 sum=00000110
* bcd_in1=01111001 bcd_in2=00101000 cout=1 sum=00000111
* bcd_in1=01111001 bcd_in2=00101001 cout=1 sum=00001000
* bcd_in1=01111001 bcd_in2=00110000 cout=1 sum=00001001
* bcd_in1=01111001 bcd_in2=00110001 cout=1 sum=00010000
* bcd_in1=01111001 bcd_in2=00110010 cout=1 sum=00010001
* bcd_in1=01111001 bcd_in2=00110011 cout=1 sum=00010010
* bcd_in1=01111001 bcd_in2=00110100 cout=1 sum=00010011
* bcd_in1=01111001 bcd_in2=00110101 cout=1 sum=00010100
* bcd_in1=01111001 bcd_in2=00110110 cout=1 sum=00010101
* bcd_in1=01111001 bcd_in2=00110111 cout=1 sum=00010110
* bcd_in1=01111001 bcd_in2=00111000 cout=1 sum=00010111
* bcd_in1=01111001 bcd_in2=00111001 cout=1 sum=00011000
* bcd_in1=01111001 bcd_in2=01000000 cout=1 sum=00011001
* bcd_in1=01111001 bcd_in2=01000001 cout=1 sum=00100000
* bcd_in1=01111001 bcd_in2=01000010 cout=1 sum=00100001
* bcd_in1=01111001 bcd_in2=01000011 cout=1 sum=00100010
* bcd_in1=01111001 bcd_in2=01000100 cout=1 sum=00100011
* bcd_in1=01111001 bcd_in2=01000101 cout=1 sum=00100100
* bcd_in1=01111001 bcd_in2=01000110 cout=1 sum=00100101
* bcd_in1=01111001 bcd_in2=01000111 cout=1 sum=00100110
* bcd_in1=01111001 bcd_in2=01001000 cout=1 sum=00100111
* bcd_in1=01111001 bcd_in2=01001001 cout=1 sum=00101000
* bcd_in1=01111001 bcd_in2=01010000 cout=1 sum=00101001
* bcd_in1=01111001 bcd_in2=01010001 cout=1 sum=00110000
* bcd_in1=01111001 bcd_in2=01010010 cout=1 sum=00110001
* bcd_in1=01111001 bcd_in2=01010011 cout=1 sum=00110010
* bcd_in1=01111001 bcd_in2=01010100 cout=1 sum=00110011
* bcd_in1=01111001 bcd_in2=01010101 cout=1 sum=00110100
* bcd_in1=01111001 bcd_in2=01010110 cout=1 sum=00110101
* bcd_in1=01111001 bcd_in2=01010111 cout=1 sum=00110110
* bcd_in1=01111001 bcd_in2=01011000 cout=1 sum=00110111
* bcd_in1=01111001 bcd_in2=01011001 cout=1 sum=00111000
* bcd_in1=01111001 bcd_in2=01100000 cout=1 sum=00111001
* bcd_in1=01111001 bcd_in2=01100001 cout=1 sum=01000000
* bcd_in1=01111001 bcd_in2=01100010 cout=1 sum=01000001
* bcd_in1=01111001 bcd_in2=01100011 cout=1 sum=01000010
* bcd_in1=01111001 bcd_in2=01100100 cout=1 sum=01000011
* bcd_in1=01111001 bcd_in2=01100101 cout=1 sum=01000100
* bcd_in1=01111001 bcd_in2=01100110 cout=1 sum=01000101
* bcd_in1=01111001 bcd_in2=01100111 cout=1 sum=01000110
* bcd_in1=01111001 bcd_in2=01101000 cout=1 sum=01000111
* bcd_in1=01111001 bcd_in2=01101001 cout=1 sum=01001000
* bcd_in1=01111001 bcd_in2=01110000 cout=1 sum=01001001
* bcd_in1=01111001 bcd_in2=01110001 cout=1 sum=01010000
* bcd_in1=01111001 bcd_in2=01110010 cout=1 sum=01010001
* bcd_in1=01111001 bcd_in2=01110011 cout=1 sum=01010010
* bcd_in1=01111001 bcd_in2=01110100 cout=1 sum=01010011
* bcd_in1=01111001 bcd_in2=01110101 cout=1 sum=01010100
* bcd_in1=01111001 bcd_in2=01110110 cout=1 sum=01010101
* bcd_in1=01111001 bcd_in2=01110111 cout=1 sum=01010110
* bcd_in1=01111001 bcd_in2=01111000 cout=1 sum=01010111
* bcd_in1=01111001 bcd_in2=01111001 cout=1 sum=01011000
* bcd_in1=01111001 bcd_in2=10000000 cout=1 sum=01011001
* bcd_in1=01111001 bcd_in2=10000001 cout=1 sum=01100000
* bcd_in1=01111001 bcd_in2=10000010 cout=1 sum=01100001
* bcd_in1=01111001 bcd_in2=10000011 cout=1 sum=01100010
* bcd_in1=01111001 bcd_in2=10000100 cout=1 sum=01100011
* bcd_in1=01111001 bcd_in2=10000101 cout=1 sum=01100100
* bcd_in1=01111001 bcd_in2=10000110 cout=1 sum=01100101
* bcd_in1=01111001 bcd_in2=10000111 cout=1 sum=01100110
* bcd_in1=01111001 bcd_in2=10001000 cout=1 sum=01100111
* bcd_in1=01111001 bcd_in2=10001001 cout=1 sum=01101000
* bcd_in1=01111001 bcd_in2=10010000 cout=1 sum=01101001
* bcd_in1=01111001 bcd_in2=10010001 cout=1 sum=01110000
* bcd_in1=01111001 bcd_in2=10010010 cout=1 sum=01110001
* bcd_in1=01111001 bcd_in2=10010011 cout=1 sum=01110010
* bcd_in1=01111001 bcd_in2=10010100 cout=1 sum=01110011
* bcd_in1=01111001 bcd_in2=10010101 cout=1 sum=01110100
* bcd_in1=01111001 bcd_in2=10010110 cout=1 sum=01110101
* bcd_in1=01111001 bcd_in2=10010111 cout=1 sum=01110110
* bcd_in1=01111001 bcd_in2=10011000 cout=1 sum=01110111
* bcd_in1=01111001 bcd_in2=10011001 cout=1 sum=01111000
* bcd_in1=10000000 bcd_in2=00000000 cout=0 sum=10000000
* bcd_in1=10000000 bcd_in2=00000001 cout=0 sum=10000001
* bcd_in1=10000000 bcd_in2=00000010 cout=0 sum=10000010
* bcd_in1=10000000 bcd_in2=00000011 cout=0 sum=10000011
* bcd_in1=10000000 bcd_in2=00000100 cout=0 sum=10000100
* bcd_in1=10000000 bcd_in2=00000101 cout=0 sum=10000101
* bcd_in1=10000000 bcd_in2=00000110 cout=0 sum=10000110
* bcd_in1=10000000 bcd_in2=00000111 cout=0 sum=10000111
* bcd_in1=10000000 bcd_in2=00001000 cout=0 sum=10001000
* bcd_in1=10000000 bcd_in2=00001001 cout=0 sum=10001001
* bcd_in1=10000000 bcd_in2=00010000 cout=0 sum=10010000
* bcd_in1=10000000 bcd_in2=00010001 cout=0 sum=10010001
* bcd_in1=10000000 bcd_in2=00010010 cout=0 sum=10010010
* bcd_in1=10000000 bcd_in2=00010011 cout=0 sum=10010011
* bcd_in1=10000000 bcd_in2=00010100 cout=0 sum=10010100
* bcd_in1=10000000 bcd_in2=00010101 cout=0 sum=10010101
* bcd_in1=10000000 bcd_in2=00010110 cout=0 sum=10010110
* bcd_in1=10000000 bcd_in2=00010111 cout=0 sum=10010111
* bcd_in1=10000000 bcd_in2=00011000 cout=0 sum=10011000
* bcd_in1=10000000 bcd_in2=00011001 cout=0 sum=10011001
* bcd_in1=10000000 bcd_in2=00100000 cout=1 sum=00000000
* bcd_in1=10000000 bcd_in2=00100001 cout=1 sum=00000001
* bcd_in1=10000000 bcd_in2=00100010 cout=1 sum=00000010
* bcd_in1=10000000 bcd_in2=00100011 cout=1 sum=00000011
* bcd_in1=10000000 bcd_in2=00100100 cout=1 sum=00000100
* bcd_in1=10000000 bcd_in2=00100101 cout=1 sum=00000101
* bcd_in1=10000000 bcd_in2=00100110 cout=1 sum=00000110
* bcd_in1=10000000 bcd_in2=00100111 cout=1 sum=00000111
* bcd_in1=10000000 bcd_in2=00101000 cout=1 sum=00001000
* bcd_in1=10000000 bcd_in2=00101001 cout=1 sum=00001001
* bcd_in1=10000000 bcd_in2=00110000 cout=1 sum=00010000
* bcd_in1=10000000 bcd_in2=00110001 cout=1 sum=00010001
* bcd_in1=10000000 bcd_in2=00110010 cout=1 sum=00010010
* bcd_in1=10000000 bcd_in2=00110011 cout=1 sum=00010011
* bcd_in1=10000000 bcd_in2=00110100 cout=1 sum=00010100
* bcd_in1=10000000 bcd_in2=00110101 cout=1 sum=00010101
* bcd_in1=10000000 bcd_in2=00110110 cout=1 sum=00010110
* bcd_in1=10000000 bcd_in2=00110111 cout=1 sum=00010111
* bcd_in1=10000000 bcd_in2=00111000 cout=1 sum=00011000
* bcd_in1=10000000 bcd_in2=00111001 cout=1 sum=00011001
* bcd_in1=10000000 bcd_in2=01000000 cout=1 sum=00100000
* bcd_in1=10000000 bcd_in2=01000001 cout=1 sum=00100001
* bcd_in1=10000000 bcd_in2=01000010 cout=1 sum=00100010
* bcd_in1=10000000 bcd_in2=01000011 cout=1 sum=00100011
* bcd_in1=10000000 bcd_in2=01000100 cout=1 sum=00100100
* bcd_in1=10000000 bcd_in2=01000101 cout=1 sum=00100101
* bcd_in1=10000000 bcd_in2=01000110 cout=1 sum=00100110
* bcd_in1=10000000 bcd_in2=01000111 cout=1 sum=00100111
* bcd_in1=10000000 bcd_in2=01001000 cout=1 sum=00101000
* bcd_in1=10000000 bcd_in2=01001001 cout=1 sum=00101001
* bcd_in1=10000000 bcd_in2=01010000 cout=1 sum=00110000
* bcd_in1=10000000 bcd_in2=01010001 cout=1 sum=00110001
* bcd_in1=10000000 bcd_in2=01010010 cout=1 sum=00110010
* bcd_in1=10000000 bcd_in2=01010011 cout=1 sum=00110011
* bcd_in1=10000000 bcd_in2=01010100 cout=1 sum=00110100
* bcd_in1=10000000 bcd_in2=01010101 cout=1 sum=00110101
* bcd_in1=10000000 bcd_in2=01010110 cout=1 sum=00110110
* bcd_in1=10000000 bcd_in2=01010111 cout=1 sum=00110111
* bcd_in1=10000000 bcd_in2=01011000 cout=1 sum=00111000
* bcd_in1=10000000 bcd_in2=01011001 cout=1 sum=00111001
* bcd_in1=10000000 bcd_in2=01100000 cout=1 sum=01000000
* bcd_in1=10000000 bcd_in2=01100001 cout=1 sum=01000001
* bcd_in1=10000000 bcd_in2=01100010 cout=1 sum=01000010
* bcd_in1=10000000 bcd_in2=01100011 cout=1 sum=01000011
* bcd_in1=10000000 bcd_in2=01100100 cout=1 sum=01000100
* bcd_in1=10000000 bcd_in2=01100101 cout=1 sum=01000101
* bcd_in1=10000000 bcd_in2=01100110 cout=1 sum=01000110
* bcd_in1=10000000 bcd_in2=01100111 cout=1 sum=01000111
* bcd_in1=10000000 bcd_in2=01101000 cout=1 sum=01001000
* bcd_in1=10000000 bcd_in2=01101001 cout=1 sum=01001001
* bcd_in1=10000000 bcd_in2=01110000 cout=1 sum=01010000
* bcd_in1=10000000 bcd_in2=01110001 cout=1 sum=01010001
* bcd_in1=10000000 bcd_in2=01110010 cout=1 sum=01010010
* bcd_in1=10000000 bcd_in2=01110011 cout=1 sum=01010011
* bcd_in1=10000000 bcd_in2=01110100 cout=1 sum=01010100
* bcd_in1=10000000 bcd_in2=01110101 cout=1 sum=01010101
* bcd_in1=10000000 bcd_in2=01110110 cout=1 sum=01010110
* bcd_in1=10000000 bcd_in2=01110111 cout=1 sum=01010111
* bcd_in1=10000000 bcd_in2=01111000 cout=1 sum=01011000
* bcd_in1=10000000 bcd_in2=01111001 cout=1 sum=01011001
* bcd_in1=10000000 bcd_in2=10000000 cout=1 sum=01100000
* bcd_in1=10000000 bcd_in2=10000001 cout=1 sum=01100001
* bcd_in1=10000000 bcd_in2=10000010 cout=1 sum=01100010
* bcd_in1=10000000 bcd_in2=10000011 cout=1 sum=01100011
* bcd_in1=10000000 bcd_in2=10000100 cout=1 sum=01100100
* bcd_in1=10000000 bcd_in2=10000101 cout=1 sum=01100101
* bcd_in1=10000000 bcd_in2=10000110 cout=1 sum=01100110
* bcd_in1=10000000 bcd_in2=10000111 cout=1 sum=01100111
* bcd_in1=10000000 bcd_in2=10001000 cout=1 sum=01101000
* bcd_in1=10000000 bcd_in2=10001001 cout=1 sum=01101001
* bcd_in1=10000000 bcd_in2=10010000 cout=1 sum=01110000
* bcd_in1=10000000 bcd_in2=10010001 cout=1 sum=01110001
* bcd_in1=10000000 bcd_in2=10010010 cout=1 sum=01110010
* bcd_in1=10000000 bcd_in2=10010011 cout=1 sum=01110011
* bcd_in1=10000000 bcd_in2=10010100 cout=1 sum=01110100
* bcd_in1=10000000 bcd_in2=10010101 cout=1 sum=01110101
* bcd_in1=10000000 bcd_in2=10010110 cout=1 sum=01110110
* bcd_in1=10000000 bcd_in2=10010111 cout=1 sum=01110111
* bcd_in1=10000000 bcd_in2=10011000 cout=1 sum=01111000
* bcd_in1=10000000 bcd_in2=10011001 cout=1 sum=01111001
* bcd_in1=10000001 bcd_in2=00000000 cout=0 sum=10000001
* bcd_in1=10000001 bcd_in2=00000001 cout=0 sum=10000010
* bcd_in1=10000001 bcd_in2=00000010 cout=0 sum=10000011
* bcd_in1=10000001 bcd_in2=00000011 cout=0 sum=10000100
* bcd_in1=10000001 bcd_in2=00000100 cout=0 sum=10000101
* bcd_in1=10000001 bcd_in2=00000101 cout=0 sum=10000110
* bcd_in1=10000001 bcd_in2=00000110 cout=0 sum=10000111
* bcd_in1=10000001 bcd_in2=00000111 cout=0 sum=10001000
* bcd_in1=10000001 bcd_in2=00001000 cout=0 sum=10001001
* bcd_in1=10000001 bcd_in2=00001001 cout=0 sum=10010000
* bcd_in1=10000001 bcd_in2=00010000 cout=0 sum=10010001
* bcd_in1=10000001 bcd_in2=00010001 cout=0 sum=10010010
* bcd_in1=10000001 bcd_in2=00010010 cout=0 sum=10010011
* bcd_in1=10000001 bcd_in2=00010011 cout=0 sum=10010100
* bcd_in1=10000001 bcd_in2=00010100 cout=0 sum=10010101
* bcd_in1=10000001 bcd_in2=00010101 cout=0 sum=10010110
* bcd_in1=10000001 bcd_in2=00010110 cout=0 sum=10010111
* bcd_in1=10000001 bcd_in2=00010111 cout=0 sum=10011000
* bcd_in1=10000001 bcd_in2=00011000 cout=0 sum=10011001
* bcd_in1=10000001 bcd_in2=00011001 cout=1 sum=00000000
* bcd_in1=10000001 bcd_in2=00100000 cout=1 sum=00000001
* bcd_in1=10000001 bcd_in2=00100001 cout=1 sum=00000010
* bcd_in1=10000001 bcd_in2=00100010 cout=1 sum=00000011
* bcd_in1=10000001 bcd_in2=00100011 cout=1 sum=00000100
* bcd_in1=10000001 bcd_in2=00100100 cout=1 sum=00000101
* bcd_in1=10000001 bcd_in2=00100101 cout=1 sum=00000110
* bcd_in1=10000001 bcd_in2=00100110 cout=1 sum=00000111
* bcd_in1=10000001 bcd_in2=00100111 cout=1 sum=00001000
* bcd_in1=10000001 bcd_in2=00101000 cout=1 sum=00001001
* bcd_in1=10000001 bcd_in2=00101001 cout=1 sum=00010000
* bcd_in1=10000001 bcd_in2=00110000 cout=1 sum=00010001
* bcd_in1=10000001 bcd_in2=00110001 cout=1 sum=00010010
* bcd_in1=10000001 bcd_in2=00110010 cout=1 sum=00010011
* bcd_in1=10000001 bcd_in2=00110011 cout=1 sum=00010100
* bcd_in1=10000001 bcd_in2=00110100 cout=1 sum=00010101
* bcd_in1=10000001 bcd_in2=00110101 cout=1 sum=00010110
* bcd_in1=10000001 bcd_in2=00110110 cout=1 sum=00010111
* bcd_in1=10000001 bcd_in2=00110111 cout=1 sum=00011000
* bcd_in1=10000001 bcd_in2=00111000 cout=1 sum=00011001
* bcd_in1=10000001 bcd_in2=00111001 cout=1 sum=00100000
* bcd_in1=10000001 bcd_in2=01000000 cout=1 sum=00100001
* bcd_in1=10000001 bcd_in2=01000001 cout=1 sum=00100010
* bcd_in1=10000001 bcd_in2=01000010 cout=1 sum=00100011
* bcd_in1=10000001 bcd_in2=01000011 cout=1 sum=00100100
* bcd_in1=10000001 bcd_in2=01000100 cout=1 sum=00100101
* bcd_in1=10000001 bcd_in2=01000101 cout=1 sum=00100110
* bcd_in1=10000001 bcd_in2=01000110 cout=1 sum=00100111
* bcd_in1=10000001 bcd_in2=01000111 cout=1 sum=00101000
* bcd_in1=10000001 bcd_in2=01001000 cout=1 sum=00101001
* bcd_in1=10000001 bcd_in2=01001001 cout=1 sum=00110000
* bcd_in1=10000001 bcd_in2=01010000 cout=1 sum=00110001
* bcd_in1=10000001 bcd_in2=01010001 cout=1 sum=00110010
* bcd_in1=10000001 bcd_in2=01010010 cout=1 sum=00110011
* bcd_in1=10000001 bcd_in2=01010011 cout=1 sum=00110100
* bcd_in1=10000001 bcd_in2=01010100 cout=1 sum=00110101
* bcd_in1=10000001 bcd_in2=01010101 cout=1 sum=00110110
* bcd_in1=10000001 bcd_in2=01010110 cout=1 sum=00110111
* bcd_in1=10000001 bcd_in2=01010111 cout=1 sum=00111000
* bcd_in1=10000001 bcd_in2=01011000 cout=1 sum=00111001
* bcd_in1=10000001 bcd_in2=01011001 cout=1 sum=01000000
* bcd_in1=10000001 bcd_in2=01100000 cout=1 sum=01000001
* bcd_in1=10000001 bcd_in2=01100001 cout=1 sum=01000010
* bcd_in1=10000001 bcd_in2=01100010 cout=1 sum=01000011
* bcd_in1=10000001 bcd_in2=01100011 cout=1 sum=01000100
* bcd_in1=10000001 bcd_in2=01100100 cout=1 sum=01000101
* bcd_in1=10000001 bcd_in2=01100101 cout=1 sum=01000110
* bcd_in1=10000001 bcd_in2=01100110 cout=1 sum=01000111
* bcd_in1=10000001 bcd_in2=01100111 cout=1 sum=01001000
* bcd_in1=10000001 bcd_in2=01101000 cout=1 sum=01001001
* bcd_in1=10000001 bcd_in2=01101001 cout=1 sum=01010000
* bcd_in1=10000001 bcd_in2=01110000 cout=1 sum=01010001
* bcd_in1=10000001 bcd_in2=01110001 cout=1 sum=01010010
* bcd_in1=10000001 bcd_in2=01110010 cout=1 sum=01010011
* bcd_in1=10000001 bcd_in2=01110011 cout=1 sum=01010100
* bcd_in1=10000001 bcd_in2=01110100 cout=1 sum=01010101
* bcd_in1=10000001 bcd_in2=01110101 cout=1 sum=01010110
* bcd_in1=10000001 bcd_in2=01110110 cout=1 sum=01010111
* bcd_in1=10000001 bcd_in2=01110111 cout=1 sum=01011000
* bcd_in1=10000001 bcd_in2=01111000 cout=1 sum=01011001
* bcd_in1=10000001 bcd_in2=01111001 cout=1 sum=01100000
* bcd_in1=10000001 bcd_in2=10000000 cout=1 sum=01100001
* bcd_in1=10000001 bcd_in2=10000001 cout=1 sum=01100010
* bcd_in1=10000001 bcd_in2=10000010 cout=1 sum=01100011
* bcd_in1=10000001 bcd_in2=10000011 cout=1 sum=01100100
* bcd_in1=10000001 bcd_in2=10000100 cout=1 sum=01100101
* bcd_in1=10000001 bcd_in2=10000101 cout=1 sum=01100110
* bcd_in1=10000001 bcd_in2=10000110 cout=1 sum=01100111
* bcd_in1=10000001 bcd_in2=10000111 cout=1 sum=01101000
* bcd_in1=10000001 bcd_in2=10001000 cout=1 sum=01101001
* bcd_in1=10000001 bcd_in2=10001001 cout=1 sum=01110000
* bcd_in1=10000001 bcd_in2=10010000 cout=1 sum=01110001
* bcd_in1=10000001 bcd_in2=10010001 cout=1 sum=01110010
* bcd_in1=10000001 bcd_in2=10010010 cout=1 sum=01110011
* bcd_in1=10000001 bcd_in2=10010011 cout=1 sum=01110100
* bcd_in1=10000001 bcd_in2=10010100 cout=1 sum=01110101
* bcd_in1=10000001 bcd_in2=10010101 cout=1 sum=01110110
* bcd_in1=10000001 bcd_in2=10010110 cout=1 sum=01110111
* bcd_in1=10000001 bcd_in2=10010111 cout=1 sum=01111000
* bcd_in1=10000001 bcd_in2=10011000 cout=1 sum=01111001
* bcd_in1=10000001 bcd_in2=10011001 cout=1 sum=10000000
* bcd_in1=10000010 bcd_in2=00000000 cout=0 sum=10000010
* bcd_in1=10000010 bcd_in2=00000001 cout=0 sum=10000011
* bcd_in1=10000010 bcd_in2=00000010 cout=0 sum=10000100
* bcd_in1=10000010 bcd_in2=00000011 cout=0 sum=10000101
* bcd_in1=10000010 bcd_in2=00000100 cout=0 sum=10000110
* bcd_in1=10000010 bcd_in2=00000101 cout=0 sum=10000111
* bcd_in1=10000010 bcd_in2=00000110 cout=0 sum=10001000
* bcd_in1=10000010 bcd_in2=00000111 cout=0 sum=10001001
* bcd_in1=10000010 bcd_in2=00001000 cout=0 sum=10010000
* bcd_in1=10000010 bcd_in2=00001001 cout=0 sum=10010001
* bcd_in1=10000010 bcd_in2=00010000 cout=0 sum=10010010
* bcd_in1=10000010 bcd_in2=00010001 cout=0 sum=10010011
* bcd_in1=10000010 bcd_in2=00010010 cout=0 sum=10010100
* bcd_in1=10000010 bcd_in2=00010011 cout=0 sum=10010101
* bcd_in1=10000010 bcd_in2=00010100 cout=0 sum=10010110
* bcd_in1=10000010 bcd_in2=00010101 cout=0 sum=10010111
* bcd_in1=10000010 bcd_in2=00010110 cout=0 sum=10011000
* bcd_in1=10000010 bcd_in2=00010111 cout=0 sum=10011001
* bcd_in1=10000010 bcd_in2=00011000 cout=1 sum=00000000
* bcd_in1=10000010 bcd_in2=00011001 cout=1 sum=00000001
* bcd_in1=10000010 bcd_in2=00100000 cout=1 sum=00000010
* bcd_in1=10000010 bcd_in2=00100001 cout=1 sum=00000011
* bcd_in1=10000010 bcd_in2=00100010 cout=1 sum=00000100
* bcd_in1=10000010 bcd_in2=00100011 cout=1 sum=00000101
* bcd_in1=10000010 bcd_in2=00100100 cout=1 sum=00000110
* bcd_in1=10000010 bcd_in2=00100101 cout=1 sum=00000111
* bcd_in1=10000010 bcd_in2=00100110 cout=1 sum=00001000
* bcd_in1=10000010 bcd_in2=00100111 cout=1 sum=00001001
* bcd_in1=10000010 bcd_in2=00101000 cout=1 sum=00010000
* bcd_in1=10000010 bcd_in2=00101001 cout=1 sum=00010001
* bcd_in1=10000010 bcd_in2=00110000 cout=1 sum=00010010
* bcd_in1=10000010 bcd_in2=00110001 cout=1 sum=00010011
* bcd_in1=10000010 bcd_in2=00110010 cout=1 sum=00010100
* bcd_in1=10000010 bcd_in2=00110011 cout=1 sum=00010101
* bcd_in1=10000010 bcd_in2=00110100 cout=1 sum=00010110
* bcd_in1=10000010 bcd_in2=00110101 cout=1 sum=00010111
* bcd_in1=10000010 bcd_in2=00110110 cout=1 sum=00011000
* bcd_in1=10000010 bcd_in2=00110111 cout=1 sum=00011001
* bcd_in1=10000010 bcd_in2=00111000 cout=1 sum=00100000
* bcd_in1=10000010 bcd_in2=00111001 cout=1 sum=00100001
* bcd_in1=10000010 bcd_in2=01000000 cout=1 sum=00100010
* bcd_in1=10000010 bcd_in2=01000001 cout=1 sum=00100011
* bcd_in1=10000010 bcd_in2=01000010 cout=1 sum=00100100
* bcd_in1=10000010 bcd_in2=01000011 cout=1 sum=00100101
* bcd_in1=10000010 bcd_in2=01000100 cout=1 sum=00100110
* bcd_in1=10000010 bcd_in2=01000101 cout=1 sum=00100111
* bcd_in1=10000010 bcd_in2=01000110 cout=1 sum=00101000
* bcd_in1=10000010 bcd_in2=01000111 cout=1 sum=00101001
* bcd_in1=10000010 bcd_in2=01001000 cout=1 sum=00110000
* bcd_in1=10000010 bcd_in2=01001001 cout=1 sum=00110001
* bcd_in1=10000010 bcd_in2=01010000 cout=1 sum=00110010
* bcd_in1=10000010 bcd_in2=01010001 cout=1 sum=00110011
* bcd_in1=10000010 bcd_in2=01010010 cout=1 sum=00110100
* bcd_in1=10000010 bcd_in2=01010011 cout=1 sum=00110101
* bcd_in1=10000010 bcd_in2=01010100 cout=1 sum=00110110
* bcd_in1=10000010 bcd_in2=01010101 cout=1 sum=00110111
* bcd_in1=10000010 bcd_in2=01010110 cout=1 sum=00111000
* bcd_in1=10000010 bcd_in2=01010111 cout=1 sum=00111001
* bcd_in1=10000010 bcd_in2=01011000 cout=1 sum=01000000
* bcd_in1=10000010 bcd_in2=01011001 cout=1 sum=01000001
* bcd_in1=10000010 bcd_in2=01100000 cout=1 sum=01000010
* bcd_in1=10000010 bcd_in2=01100001 cout=1 sum=01000011
* bcd_in1=10000010 bcd_in2=01100010 cout=1 sum=01000100
* bcd_in1=10000010 bcd_in2=01100011 cout=1 sum=01000101
* bcd_in1=10000010 bcd_in2=01100100 cout=1 sum=01000110
* bcd_in1=10000010 bcd_in2=01100101 cout=1 sum=01000111
* bcd_in1=10000010 bcd_in2=01100110 cout=1 sum=01001000
* bcd_in1=10000010 bcd_in2=01100111 cout=1 sum=01001001
* bcd_in1=10000010 bcd_in2=01101000 cout=1 sum=01010000
* bcd_in1=10000010 bcd_in2=01101001 cout=1 sum=01010001
* bcd_in1=10000010 bcd_in2=01110000 cout=1 sum=01010010
* bcd_in1=10000010 bcd_in2=01110001 cout=1 sum=01010011
* bcd_in1=10000010 bcd_in2=01110010 cout=1 sum=01010100
* bcd_in1=10000010 bcd_in2=01110011 cout=1 sum=01010101
* bcd_in1=10000010 bcd_in2=01110100 cout=1 sum=01010110
* bcd_in1=10000010 bcd_in2=01110101 cout=1 sum=01010111
* bcd_in1=10000010 bcd_in2=01110110 cout=1 sum=01011000
* bcd_in1=10000010 bcd_in2=01110111 cout=1 sum=01011001
* bcd_in1=10000010 bcd_in2=01111000 cout=1 sum=01100000
* bcd_in1=10000010 bcd_in2=01111001 cout=1 sum=01100001
* bcd_in1=10000010 bcd_in2=10000000 cout=1 sum=01100010
* bcd_in1=10000010 bcd_in2=10000001 cout=1 sum=01100011
* bcd_in1=10000010 bcd_in2=10000010 cout=1 sum=01100100
* bcd_in1=10000010 bcd_in2=10000011 cout=1 sum=01100101
* bcd_in1=10000010 bcd_in2=10000100 cout=1 sum=01100110
* bcd_in1=10000010 bcd_in2=10000101 cout=1 sum=01100111
* bcd_in1=10000010 bcd_in2=10000110 cout=1 sum=01101000
* bcd_in1=10000010 bcd_in2=10000111 cout=1 sum=01101001
* bcd_in1=10000010 bcd_in2=10001000 cout=1 sum=01110000
* bcd_in1=10000010 bcd_in2=10001001 cout=1 sum=01110001
* bcd_in1=10000010 bcd_in2=10010000 cout=1 sum=01110010
* bcd_in1=10000010 bcd_in2=10010001 cout=1 sum=01110011
* bcd_in1=10000010 bcd_in2=10010010 cout=1 sum=01110100
* bcd_in1=10000010 bcd_in2=10010011 cout=1 sum=01110101
* bcd_in1=10000010 bcd_in2=10010100 cout=1 sum=01110110
* bcd_in1=10000010 bcd_in2=10010101 cout=1 sum=01110111
* bcd_in1=10000010 bcd_in2=10010110 cout=1 sum=01111000
* bcd_in1=10000010 bcd_in2=10010111 cout=1 sum=01111001
* bcd_in1=10000010 bcd_in2=10011000 cout=1 sum=10000000
* bcd_in1=10000010 bcd_in2=10011001 cout=1 sum=10000001
* bcd_in1=10000011 bcd_in2=00000000 cout=0 sum=10000011
* bcd_in1=10000011 bcd_in2=00000001 cout=0 sum=10000100
* bcd_in1=10000011 bcd_in2=00000010 cout=0 sum=10000101
* bcd_in1=10000011 bcd_in2=00000011 cout=0 sum=10000110
* bcd_in1=10000011 bcd_in2=00000100 cout=0 sum=10000111
* bcd_in1=10000011 bcd_in2=00000101 cout=0 sum=10001000
* bcd_in1=10000011 bcd_in2=00000110 cout=0 sum=10001001
* bcd_in1=10000011 bcd_in2=00000111 cout=0 sum=10010000
* bcd_in1=10000011 bcd_in2=00001000 cout=0 sum=10010001
* bcd_in1=10000011 bcd_in2=00001001 cout=0 sum=10010010
* bcd_in1=10000011 bcd_in2=00010000 cout=0 sum=10010011
* bcd_in1=10000011 bcd_in2=00010001 cout=0 sum=10010100
* bcd_in1=10000011 bcd_in2=00010010 cout=0 sum=10010101
* bcd_in1=10000011 bcd_in2=00010011 cout=0 sum=10010110
* bcd_in1=10000011 bcd_in2=00010100 cout=0 sum=10010111
* bcd_in1=10000011 bcd_in2=00010101 cout=0 sum=10011000
* bcd_in1=10000011 bcd_in2=00010110 cout=0 sum=10011001
* bcd_in1=10000011 bcd_in2=00010111 cout=1 sum=00000000
* bcd_in1=10000011 bcd_in2=00011000 cout=1 sum=00000001
* bcd_in1=10000011 bcd_in2=00011001 cout=1 sum=00000010
* bcd_in1=10000011 bcd_in2=00100000 cout=1 sum=00000011
* bcd_in1=10000011 bcd_in2=00100001 cout=1 sum=00000100
* bcd_in1=10000011 bcd_in2=00100010 cout=1 sum=00000101
* bcd_in1=10000011 bcd_in2=00100011 cout=1 sum=00000110
* bcd_in1=10000011 bcd_in2=00100100 cout=1 sum=00000111
* bcd_in1=10000011 bcd_in2=00100101 cout=1 sum=00001000
* bcd_in1=10000011 bcd_in2=00100110 cout=1 sum=00001001
* bcd_in1=10000011 bcd_in2=00100111 cout=1 sum=00010000
* bcd_in1=10000011 bcd_in2=00101000 cout=1 sum=00010001
* bcd_in1=10000011 bcd_in2=00101001 cout=1 sum=00010010
* bcd_in1=10000011 bcd_in2=00110000 cout=1 sum=00010011
* bcd_in1=10000011 bcd_in2=00110001 cout=1 sum=00010100
* bcd_in1=10000011 bcd_in2=00110010 cout=1 sum=00010101
* bcd_in1=10000011 bcd_in2=00110011 cout=1 sum=00010110
* bcd_in1=10000011 bcd_in2=00110100 cout=1 sum=00010111
* bcd_in1=10000011 bcd_in2=00110101 cout=1 sum=00011000
* bcd_in1=10000011 bcd_in2=00110110 cout=1 sum=00011001
* bcd_in1=10000011 bcd_in2=00110111 cout=1 sum=00100000
* bcd_in1=10000011 bcd_in2=00111000 cout=1 sum=00100001
* bcd_in1=10000011 bcd_in2=00111001 cout=1 sum=00100010
* bcd_in1=10000011 bcd_in2=01000000 cout=1 sum=00100011
* bcd_in1=10000011 bcd_in2=01000001 cout=1 sum=00100100
* bcd_in1=10000011 bcd_in2=01000010 cout=1 sum=00100101
* bcd_in1=10000011 bcd_in2=01000011 cout=1 sum=00100110
* bcd_in1=10000011 bcd_in2=01000100 cout=1 sum=00100111
* bcd_in1=10000011 bcd_in2=01000101 cout=1 sum=00101000
* bcd_in1=10000011 bcd_in2=01000110 cout=1 sum=00101001
* bcd_in1=10000011 bcd_in2=01000111 cout=1 sum=00110000
* bcd_in1=10000011 bcd_in2=01001000 cout=1 sum=00110001
* bcd_in1=10000011 bcd_in2=01001001 cout=1 sum=00110010
* bcd_in1=10000011 bcd_in2=01010000 cout=1 sum=00110011
* bcd_in1=10000011 bcd_in2=01010001 cout=1 sum=00110100
* bcd_in1=10000011 bcd_in2=01010010 cout=1 sum=00110101
* bcd_in1=10000011 bcd_in2=01010011 cout=1 sum=00110110
* bcd_in1=10000011 bcd_in2=01010100 cout=1 sum=00110111
* bcd_in1=10000011 bcd_in2=01010101 cout=1 sum=00111000
* bcd_in1=10000011 bcd_in2=01010110 cout=1 sum=00111001
* bcd_in1=10000011 bcd_in2=01010111 cout=1 sum=01000000
* bcd_in1=10000011 bcd_in2=01011000 cout=1 sum=01000001
* bcd_in1=10000011 bcd_in2=01011001 cout=1 sum=01000010
* bcd_in1=10000011 bcd_in2=01100000 cout=1 sum=01000011
* bcd_in1=10000011 bcd_in2=01100001 cout=1 sum=01000100
* bcd_in1=10000011 bcd_in2=01100010 cout=1 sum=01000101
* bcd_in1=10000011 bcd_in2=01100011 cout=1 sum=01000110
* bcd_in1=10000011 bcd_in2=01100100 cout=1 sum=01000111
* bcd_in1=10000011 bcd_in2=01100101 cout=1 sum=01001000
* bcd_in1=10000011 bcd_in2=01100110 cout=1 sum=01001001
* bcd_in1=10000011 bcd_in2=01100111 cout=1 sum=01010000
* bcd_in1=10000011 bcd_in2=01101000 cout=1 sum=01010001
* bcd_in1=10000011 bcd_in2=01101001 cout=1 sum=01010010
* bcd_in1=10000011 bcd_in2=01110000 cout=1 sum=01010011
* bcd_in1=10000011 bcd_in2=01110001 cout=1 sum=01010100
* bcd_in1=10000011 bcd_in2=01110010 cout=1 sum=01010101
* bcd_in1=10000011 bcd_in2=01110011 cout=1 sum=01010110
* bcd_in1=10000011 bcd_in2=01110100 cout=1 sum=01010111
* bcd_in1=10000011 bcd_in2=01110101 cout=1 sum=01011000
* bcd_in1=10000011 bcd_in2=01110110 cout=1 sum=01011001
* bcd_in1=10000011 bcd_in2=01110111 cout=1 sum=01100000
* bcd_in1=10000011 bcd_in2=01111000 cout=1 sum=01100001
* bcd_in1=10000011 bcd_in2=01111001 cout=1 sum=01100010
* bcd_in1=10000011 bcd_in2=10000000 cout=1 sum=01100011
* bcd_in1=10000011 bcd_in2=10000001 cout=1 sum=01100100
* bcd_in1=10000011 bcd_in2=10000010 cout=1 sum=01100101
* bcd_in1=10000011 bcd_in2=10000011 cout=1 sum=01100110
* bcd_in1=10000011 bcd_in2=10000100 cout=1 sum=01100111
* bcd_in1=10000011 bcd_in2=10000101 cout=1 sum=01101000
* bcd_in1=10000011 bcd_in2=10000110 cout=1 sum=01101001
* bcd_in1=10000011 bcd_in2=10000111 cout=1 sum=01110000
* bcd_in1=10000011 bcd_in2=10001000 cout=1 sum=01110001
* bcd_in1=10000011 bcd_in2=10001001 cout=1 sum=01110010
* bcd_in1=10000011 bcd_in2=10010000 cout=1 sum=01110011
* bcd_in1=10000011 bcd_in2=10010001 cout=1 sum=01110100
* bcd_in1=10000011 bcd_in2=10010010 cout=1 sum=01110101
* bcd_in1=10000011 bcd_in2=10010011 cout=1 sum=01110110
* bcd_in1=10000011 bcd_in2=10010100 cout=1 sum=01110111
* bcd_in1=10000011 bcd_in2=10010101 cout=1 sum=01111000
* bcd_in1=10000011 bcd_in2=10010110 cout=1 sum=01111001
* bcd_in1=10000011 bcd_in2=10010111 cout=1 sum=10000000
* bcd_in1=10000011 bcd_in2=10011000 cout=1 sum=10000001
* bcd_in1=10000011 bcd_in2=10011001 cout=1 sum=10000010
* bcd_in1=10000100 bcd_in2=00000000 cout=0 sum=10000100
* bcd_in1=10000100 bcd_in2=00000001 cout=0 sum=10000101
* bcd_in1=10000100 bcd_in2=00000010 cout=0 sum=10000110
* bcd_in1=10000100 bcd_in2=00000011 cout=0 sum=10000111
* bcd_in1=10000100 bcd_in2=00000100 cout=0 sum=10001000
* bcd_in1=10000100 bcd_in2=00000101 cout=0 sum=10001001
* bcd_in1=10000100 bcd_in2=00000110 cout=0 sum=10010000
* bcd_in1=10000100 bcd_in2=00000111 cout=0 sum=10010001
* bcd_in1=10000100 bcd_in2=00001000 cout=0 sum=10010010
* bcd_in1=10000100 bcd_in2=00001001 cout=0 sum=10010011
* bcd_in1=10000100 bcd_in2=00010000 cout=0 sum=10010100
* bcd_in1=10000100 bcd_in2=00010001 cout=0 sum=10010101
* bcd_in1=10000100 bcd_in2=00010010 cout=0 sum=10010110
* bcd_in1=10000100 bcd_in2=00010011 cout=0 sum=10010111
* bcd_in1=10000100 bcd_in2=00010100 cout=0 sum=10011000
* bcd_in1=10000100 bcd_in2=00010101 cout=0 sum=10011001
* bcd_in1=10000100 bcd_in2=00010110 cout=1 sum=00000000
* bcd_in1=10000100 bcd_in2=00010111 cout=1 sum=00000001
* bcd_in1=10000100 bcd_in2=00011000 cout=1 sum=00000010
* bcd_in1=10000100 bcd_in2=00011001 cout=1 sum=00000011
* bcd_in1=10000100 bcd_in2=00100000 cout=1 sum=00000100
* bcd_in1=10000100 bcd_in2=00100001 cout=1 sum=00000101
* bcd_in1=10000100 bcd_in2=00100010 cout=1 sum=00000110
* bcd_in1=10000100 bcd_in2=00100011 cout=1 sum=00000111
* bcd_in1=10000100 bcd_in2=00100100 cout=1 sum=00001000
* bcd_in1=10000100 bcd_in2=00100101 cout=1 sum=00001001
* bcd_in1=10000100 bcd_in2=00100110 cout=1 sum=00010000
* bcd_in1=10000100 bcd_in2=00100111 cout=1 sum=00010001
* bcd_in1=10000100 bcd_in2=00101000 cout=1 sum=00010010
* bcd_in1=10000100 bcd_in2=00101001 cout=1 sum=00010011
* bcd_in1=10000100 bcd_in2=00110000 cout=1 sum=00010100
* bcd_in1=10000100 bcd_in2=00110001 cout=1 sum=00010101
* bcd_in1=10000100 bcd_in2=00110010 cout=1 sum=00010110
* bcd_in1=10000100 bcd_in2=00110011 cout=1 sum=00010111
* bcd_in1=10000100 bcd_in2=00110100 cout=1 sum=00011000
* bcd_in1=10000100 bcd_in2=00110101 cout=1 sum=00011001
* bcd_in1=10000100 bcd_in2=00110110 cout=1 sum=00100000
* bcd_in1=10000100 bcd_in2=00110111 cout=1 sum=00100001
* bcd_in1=10000100 bcd_in2=00111000 cout=1 sum=00100010
* bcd_in1=10000100 bcd_in2=00111001 cout=1 sum=00100011
* bcd_in1=10000100 bcd_in2=01000000 cout=1 sum=00100100
* bcd_in1=10000100 bcd_in2=01000001 cout=1 sum=00100101
* bcd_in1=10000100 bcd_in2=01000010 cout=1 sum=00100110
* bcd_in1=10000100 bcd_in2=01000011 cout=1 sum=00100111
* bcd_in1=10000100 bcd_in2=01000100 cout=1 sum=00101000
* bcd_in1=10000100 bcd_in2=01000101 cout=1 sum=00101001
* bcd_in1=10000100 bcd_in2=01000110 cout=1 sum=00110000
* bcd_in1=10000100 bcd_in2=01000111 cout=1 sum=00110001
* bcd_in1=10000100 bcd_in2=01001000 cout=1 sum=00110010
* bcd_in1=10000100 bcd_in2=01001001 cout=1 sum=00110011
* bcd_in1=10000100 bcd_in2=01010000 cout=1 sum=00110100
* bcd_in1=10000100 bcd_in2=01010001 cout=1 sum=00110101
* bcd_in1=10000100 bcd_in2=01010010 cout=1 sum=00110110
* bcd_in1=10000100 bcd_in2=01010011 cout=1 sum=00110111
* bcd_in1=10000100 bcd_in2=01010100 cout=1 sum=00111000
* bcd_in1=10000100 bcd_in2=01010101 cout=1 sum=00111001
* bcd_in1=10000100 bcd_in2=01010110 cout=1 sum=01000000
* bcd_in1=10000100 bcd_in2=01010111 cout=1 sum=01000001
* bcd_in1=10000100 bcd_in2=01011000 cout=1 sum=01000010
* bcd_in1=10000100 bcd_in2=01011001 cout=1 sum=01000011
* bcd_in1=10000100 bcd_in2=01100000 cout=1 sum=01000100
* bcd_in1=10000100 bcd_in2=01100001 cout=1 sum=01000101
* bcd_in1=10000100 bcd_in2=01100010 cout=1 sum=01000110
* bcd_in1=10000100 bcd_in2=01100011 cout=1 sum=01000111
* bcd_in1=10000100 bcd_in2=01100100 cout=1 sum=01001000
* bcd_in1=10000100 bcd_in2=01100101 cout=1 sum=01001001
* bcd_in1=10000100 bcd_in2=01100110 cout=1 sum=01010000
* bcd_in1=10000100 bcd_in2=01100111 cout=1 sum=01010001
* bcd_in1=10000100 bcd_in2=01101000 cout=1 sum=01010010
* bcd_in1=10000100 bcd_in2=01101001 cout=1 sum=01010011
* bcd_in1=10000100 bcd_in2=01110000 cout=1 sum=01010100
* bcd_in1=10000100 bcd_in2=01110001 cout=1 sum=01010101
* bcd_in1=10000100 bcd_in2=01110010 cout=1 sum=01010110
* bcd_in1=10000100 bcd_in2=01110011 cout=1 sum=01010111
* bcd_in1=10000100 bcd_in2=01110100 cout=1 sum=01011000
* bcd_in1=10000100 bcd_in2=01110101 cout=1 sum=01011001
* bcd_in1=10000100 bcd_in2=01110110 cout=1 sum=01100000
* bcd_in1=10000100 bcd_in2=01110111 cout=1 sum=01100001
* bcd_in1=10000100 bcd_in2=01111000 cout=1 sum=01100010
* bcd_in1=10000100 bcd_in2=01111001 cout=1 sum=01100011
* bcd_in1=10000100 bcd_in2=10000000 cout=1 sum=01100100
* bcd_in1=10000100 bcd_in2=10000001 cout=1 sum=01100101
* bcd_in1=10000100 bcd_in2=10000010 cout=1 sum=01100110
* bcd_in1=10000100 bcd_in2=10000011 cout=1 sum=01100111
* bcd_in1=10000100 bcd_in2=10000100 cout=1 sum=01101000
* bcd_in1=10000100 bcd_in2=10000101 cout=1 sum=01101001
* bcd_in1=10000100 bcd_in2=10000110 cout=1 sum=01110000
* bcd_in1=10000100 bcd_in2=10000111 cout=1 sum=01110001
* bcd_in1=10000100 bcd_in2=10001000 cout=1 sum=01110010
* bcd_in1=10000100 bcd_in2=10001001 cout=1 sum=01110011
* bcd_in1=10000100 bcd_in2=10010000 cout=1 sum=01110100
* bcd_in1=10000100 bcd_in2=10010001 cout=1 sum=01110101
* bcd_in1=10000100 bcd_in2=10010010 cout=1 sum=01110110
* bcd_in1=10000100 bcd_in2=10010011 cout=1 sum=01110111
* bcd_in1=10000100 bcd_in2=10010100 cout=1 sum=01111000
* bcd_in1=10000100 bcd_in2=10010101 cout=1 sum=01111001
* bcd_in1=10000100 bcd_in2=10010110 cout=1 sum=10000000
* bcd_in1=10000100 bcd_in2=10010111 cout=1 sum=10000001
* bcd_in1=10000100 bcd_in2=10011000 cout=1 sum=10000010
* bcd_in1=10000100 bcd_in2=10011001 cout=1 sum=10000011
* bcd_in1=10000101 bcd_in2=00000000 cout=0 sum=10000101
* bcd_in1=10000101 bcd_in2=00000001 cout=0 sum=10000110
* bcd_in1=10000101 bcd_in2=00000010 cout=0 sum=10000111
* bcd_in1=10000101 bcd_in2=00000011 cout=0 sum=10001000
* bcd_in1=10000101 bcd_in2=00000100 cout=0 sum=10001001
* bcd_in1=10000101 bcd_in2=00000101 cout=0 sum=10010000
* bcd_in1=10000101 bcd_in2=00000110 cout=0 sum=10010001
* bcd_in1=10000101 bcd_in2=00000111 cout=0 sum=10010010
* bcd_in1=10000101 bcd_in2=00001000 cout=0 sum=10010011
* bcd_in1=10000101 bcd_in2=00001001 cout=0 sum=10010100
* bcd_in1=10000101 bcd_in2=00010000 cout=0 sum=10010101
* bcd_in1=10000101 bcd_in2=00010001 cout=0 sum=10010110
* bcd_in1=10000101 bcd_in2=00010010 cout=0 sum=10010111
* bcd_in1=10000101 bcd_in2=00010011 cout=0 sum=10011000
* bcd_in1=10000101 bcd_in2=00010100 cout=0 sum=10011001
* bcd_in1=10000101 bcd_in2=00010101 cout=1 sum=00000000
* bcd_in1=10000101 bcd_in2=00010110 cout=1 sum=00000001
* bcd_in1=10000101 bcd_in2=00010111 cout=1 sum=00000010
* bcd_in1=10000101 bcd_in2=00011000 cout=1 sum=00000011
* bcd_in1=10000101 bcd_in2=00011001 cout=1 sum=00000100
* bcd_in1=10000101 bcd_in2=00100000 cout=1 sum=00000101
* bcd_in1=10000101 bcd_in2=00100001 cout=1 sum=00000110
* bcd_in1=10000101 bcd_in2=00100010 cout=1 sum=00000111
* bcd_in1=10000101 bcd_in2=00100011 cout=1 sum=00001000
* bcd_in1=10000101 bcd_in2=00100100 cout=1 sum=00001001
* bcd_in1=10000101 bcd_in2=00100101 cout=1 sum=00010000
* bcd_in1=10000101 bcd_in2=00100110 cout=1 sum=00010001
* bcd_in1=10000101 bcd_in2=00100111 cout=1 sum=00010010
* bcd_in1=10000101 bcd_in2=00101000 cout=1 sum=00010011
* bcd_in1=10000101 bcd_in2=00101001 cout=1 sum=00010100
* bcd_in1=10000101 bcd_in2=00110000 cout=1 sum=00010101
* bcd_in1=10000101 bcd_in2=00110001 cout=1 sum=00010110
* bcd_in1=10000101 bcd_in2=00110010 cout=1 sum=00010111
* bcd_in1=10000101 bcd_in2=00110011 cout=1 sum=00011000
* bcd_in1=10000101 bcd_in2=00110100 cout=1 sum=00011001
* bcd_in1=10000101 bcd_in2=00110101 cout=1 sum=00100000
* bcd_in1=10000101 bcd_in2=00110110 cout=1 sum=00100001
* bcd_in1=10000101 bcd_in2=00110111 cout=1 sum=00100010
* bcd_in1=10000101 bcd_in2=00111000 cout=1 sum=00100011
* bcd_in1=10000101 bcd_in2=00111001 cout=1 sum=00100100
* bcd_in1=10000101 bcd_in2=01000000 cout=1 sum=00100101
* bcd_in1=10000101 bcd_in2=01000001 cout=1 sum=00100110
* bcd_in1=10000101 bcd_in2=01000010 cout=1 sum=00100111
* bcd_in1=10000101 bcd_in2=01000011 cout=1 sum=00101000
* bcd_in1=10000101 bcd_in2=01000100 cout=1 sum=00101001
* bcd_in1=10000101 bcd_in2=01000101 cout=1 sum=00110000
* bcd_in1=10000101 bcd_in2=01000110 cout=1 sum=00110001
* bcd_in1=10000101 bcd_in2=01000111 cout=1 sum=00110010
* bcd_in1=10000101 bcd_in2=01001000 cout=1 sum=00110011
* bcd_in1=10000101 bcd_in2=01001001 cout=1 sum=00110100
* bcd_in1=10000101 bcd_in2=01010000 cout=1 sum=00110101
* bcd_in1=10000101 bcd_in2=01010001 cout=1 sum=00110110
* bcd_in1=10000101 bcd_in2=01010010 cout=1 sum=00110111
* bcd_in1=10000101 bcd_in2=01010011 cout=1 sum=00111000
* bcd_in1=10000101 bcd_in2=01010100 cout=1 sum=00111001
* bcd_in1=10000101 bcd_in2=01010101 cout=1 sum=01000000
* bcd_in1=10000101 bcd_in2=01010110 cout=1 sum=01000001
* bcd_in1=10000101 bcd_in2=01010111 cout=1 sum=01000010
* bcd_in1=10000101 bcd_in2=01011000 cout=1 sum=01000011
* bcd_in1=10000101 bcd_in2=01011001 cout=1 sum=01000100
* bcd_in1=10000101 bcd_in2=01100000 cout=1 sum=01000101
* bcd_in1=10000101 bcd_in2=01100001 cout=1 sum=01000110
* bcd_in1=10000101 bcd_in2=01100010 cout=1 sum=01000111
* bcd_in1=10000101 bcd_in2=01100011 cout=1 sum=01001000
* bcd_in1=10000101 bcd_in2=01100100 cout=1 sum=01001001
* bcd_in1=10000101 bcd_in2=01100101 cout=1 sum=01010000
* bcd_in1=10000101 bcd_in2=01100110 cout=1 sum=01010001
* bcd_in1=10000101 bcd_in2=01100111 cout=1 sum=01010010
* bcd_in1=10000101 bcd_in2=01101000 cout=1 sum=01010011
* bcd_in1=10000101 bcd_in2=01101001 cout=1 sum=01010100
* bcd_in1=10000101 bcd_in2=01110000 cout=1 sum=01010101
* bcd_in1=10000101 bcd_in2=01110001 cout=1 sum=01010110
* bcd_in1=10000101 bcd_in2=01110010 cout=1 sum=01010111
* bcd_in1=10000101 bcd_in2=01110011 cout=1 sum=01011000
* bcd_in1=10000101 bcd_in2=01110100 cout=1 sum=01011001
* bcd_in1=10000101 bcd_in2=01110101 cout=1 sum=01100000
* bcd_in1=10000101 bcd_in2=01110110 cout=1 sum=01100001
* bcd_in1=10000101 bcd_in2=01110111 cout=1 sum=01100010
* bcd_in1=10000101 bcd_in2=01111000 cout=1 sum=01100011
* bcd_in1=10000101 bcd_in2=01111001 cout=1 sum=01100100
* bcd_in1=10000101 bcd_in2=10000000 cout=1 sum=01100101
* bcd_in1=10000101 bcd_in2=10000001 cout=1 sum=01100110
* bcd_in1=10000101 bcd_in2=10000010 cout=1 sum=01100111
* bcd_in1=10000101 bcd_in2=10000011 cout=1 sum=01101000
* bcd_in1=10000101 bcd_in2=10000100 cout=1 sum=01101001
* bcd_in1=10000101 bcd_in2=10000101 cout=1 sum=01110000
* bcd_in1=10000101 bcd_in2=10000110 cout=1 sum=01110001
* bcd_in1=10000101 bcd_in2=10000111 cout=1 sum=01110010
* bcd_in1=10000101 bcd_in2=10001000 cout=1 sum=01110011
* bcd_in1=10000101 bcd_in2=10001001 cout=1 sum=01110100
* bcd_in1=10000101 bcd_in2=10010000 cout=1 sum=01110101
* bcd_in1=10000101 bcd_in2=10010001 cout=1 sum=01110110
* bcd_in1=10000101 bcd_in2=10010010 cout=1 sum=01110111
* bcd_in1=10000101 bcd_in2=10010011 cout=1 sum=01111000
* bcd_in1=10000101 bcd_in2=10010100 cout=1 sum=01111001
* bcd_in1=10000101 bcd_in2=10010101 cout=1 sum=10000000
* bcd_in1=10000101 bcd_in2=10010110 cout=1 sum=10000001
* bcd_in1=10000101 bcd_in2=10010111 cout=1 sum=10000010
* bcd_in1=10000101 bcd_in2=10011000 cout=1 sum=10000011
* bcd_in1=10000101 bcd_in2=10011001 cout=1 sum=10000100
* bcd_in1=10000110 bcd_in2=00000000 cout=0 sum=10000110
* bcd_in1=10000110 bcd_in2=00000001 cout=0 sum=10000111
* bcd_in1=10000110 bcd_in2=00000010 cout=0 sum=10001000
* bcd_in1=10000110 bcd_in2=00000011 cout=0 sum=10001001
* bcd_in1=10000110 bcd_in2=00000100 cout=0 sum=10010000
* bcd_in1=10000110 bcd_in2=00000101 cout=0 sum=10010001
* bcd_in1=10000110 bcd_in2=00000110 cout=0 sum=10010010
* bcd_in1=10000110 bcd_in2=00000111 cout=0 sum=10010011
* bcd_in1=10000110 bcd_in2=00001000 cout=0 sum=10010100
* bcd_in1=10000110 bcd_in2=00001001 cout=0 sum=10010101
* bcd_in1=10000110 bcd_in2=00010000 cout=0 sum=10010110
* bcd_in1=10000110 bcd_in2=00010001 cout=0 sum=10010111
* bcd_in1=10000110 bcd_in2=00010010 cout=0 sum=10011000
* bcd_in1=10000110 bcd_in2=00010011 cout=0 sum=10011001
* bcd_in1=10000110 bcd_in2=00010100 cout=1 sum=00000000
* bcd_in1=10000110 bcd_in2=00010101 cout=1 sum=00000001
* bcd_in1=10000110 bcd_in2=00010110 cout=1 sum=00000010
* bcd_in1=10000110 bcd_in2=00010111 cout=1 sum=00000011
* bcd_in1=10000110 bcd_in2=00011000 cout=1 sum=00000100
* bcd_in1=10000110 bcd_in2=00011001 cout=1 sum=00000101
* bcd_in1=10000110 bcd_in2=00100000 cout=1 sum=00000110
* bcd_in1=10000110 bcd_in2=00100001 cout=1 sum=00000111
* bcd_in1=10000110 bcd_in2=00100010 cout=1 sum=00001000
* bcd_in1=10000110 bcd_in2=00100011 cout=1 sum=00001001
* bcd_in1=10000110 bcd_in2=00100100 cout=1 sum=00010000
* bcd_in1=10000110 bcd_in2=00100101 cout=1 sum=00010001
* bcd_in1=10000110 bcd_in2=00100110 cout=1 sum=00010010
* bcd_in1=10000110 bcd_in2=00100111 cout=1 sum=00010011
* bcd_in1=10000110 bcd_in2=00101000 cout=1 sum=00010100
* bcd_in1=10000110 bcd_in2=00101001 cout=1 sum=00010101
* bcd_in1=10000110 bcd_in2=00110000 cout=1 sum=00010110
* bcd_in1=10000110 bcd_in2=00110001 cout=1 sum=00010111
* bcd_in1=10000110 bcd_in2=00110010 cout=1 sum=00011000
* bcd_in1=10000110 bcd_in2=00110011 cout=1 sum=00011001
* bcd_in1=10000110 bcd_in2=00110100 cout=1 sum=00100000
* bcd_in1=10000110 bcd_in2=00110101 cout=1 sum=00100001
* bcd_in1=10000110 bcd_in2=00110110 cout=1 sum=00100010
* bcd_in1=10000110 bcd_in2=00110111 cout=1 sum=00100011
* bcd_in1=10000110 bcd_in2=00111000 cout=1 sum=00100100
* bcd_in1=10000110 bcd_in2=00111001 cout=1 sum=00100101
* bcd_in1=10000110 bcd_in2=01000000 cout=1 sum=00100110
* bcd_in1=10000110 bcd_in2=01000001 cout=1 sum=00100111
* bcd_in1=10000110 bcd_in2=01000010 cout=1 sum=00101000
* bcd_in1=10000110 bcd_in2=01000011 cout=1 sum=00101001
* bcd_in1=10000110 bcd_in2=01000100 cout=1 sum=00110000
* bcd_in1=10000110 bcd_in2=01000101 cout=1 sum=00110001
* bcd_in1=10000110 bcd_in2=01000110 cout=1 sum=00110010
* bcd_in1=10000110 bcd_in2=01000111 cout=1 sum=00110011
* bcd_in1=10000110 bcd_in2=01001000 cout=1 sum=00110100
* bcd_in1=10000110 bcd_in2=01001001 cout=1 sum=00110101
* bcd_in1=10000110 bcd_in2=01010000 cout=1 sum=00110110
* bcd_in1=10000110 bcd_in2=01010001 cout=1 sum=00110111
* bcd_in1=10000110 bcd_in2=01010010 cout=1 sum=00111000
* bcd_in1=10000110 bcd_in2=01010011 cout=1 sum=00111001
* bcd_in1=10000110 bcd_in2=01010100 cout=1 sum=01000000
* bcd_in1=10000110 bcd_in2=01010101 cout=1 sum=01000001
* bcd_in1=10000110 bcd_in2=01010110 cout=1 sum=01000010
* bcd_in1=10000110 bcd_in2=01010111 cout=1 sum=01000011
* bcd_in1=10000110 bcd_in2=01011000 cout=1 sum=01000100
* bcd_in1=10000110 bcd_in2=01011001 cout=1 sum=01000101
* bcd_in1=10000110 bcd_in2=01100000 cout=1 sum=01000110
* bcd_in1=10000110 bcd_in2=01100001 cout=1 sum=01000111
* bcd_in1=10000110 bcd_in2=01100010 cout=1 sum=01001000
* bcd_in1=10000110 bcd_in2=01100011 cout=1 sum=01001001
* bcd_in1=10000110 bcd_in2=01100100 cout=1 sum=01010000
* bcd_in1=10000110 bcd_in2=01100101 cout=1 sum=01010001
* bcd_in1=10000110 bcd_in2=01100110 cout=1 sum=01010010
* bcd_in1=10000110 bcd_in2=01100111 cout=1 sum=01010011
* bcd_in1=10000110 bcd_in2=01101000 cout=1 sum=01010100
* bcd_in1=10000110 bcd_in2=01101001 cout=1 sum=01010101
* bcd_in1=10000110 bcd_in2=01110000 cout=1 sum=01010110
* bcd_in1=10000110 bcd_in2=01110001 cout=1 sum=01010111
* bcd_in1=10000110 bcd_in2=01110010 cout=1 sum=01011000
* bcd_in1=10000110 bcd_in2=01110011 cout=1 sum=01011001
* bcd_in1=10000110 bcd_in2=01110100 cout=1 sum=01100000
* bcd_in1=10000110 bcd_in2=01110101 cout=1 sum=01100001
* bcd_in1=10000110 bcd_in2=01110110 cout=1 sum=01100010
* bcd_in1=10000110 bcd_in2=01110111 cout=1 sum=01100011
* bcd_in1=10000110 bcd_in2=01111000 cout=1 sum=01100100
* bcd_in1=10000110 bcd_in2=01111001 cout=1 sum=01100101
* bcd_in1=10000110 bcd_in2=10000000 cout=1 sum=01100110
* bcd_in1=10000110 bcd_in2=10000001 cout=1 sum=01100111
* bcd_in1=10000110 bcd_in2=10000010 cout=1 sum=01101000
* bcd_in1=10000110 bcd_in2=10000011 cout=1 sum=01101001
* bcd_in1=10000110 bcd_in2=10000100 cout=1 sum=01110000
* bcd_in1=10000110 bcd_in2=10000101 cout=1 sum=01110001
* bcd_in1=10000110 bcd_in2=10000110 cout=1 sum=01110010
* bcd_in1=10000110 bcd_in2=10000111 cout=1 sum=01110011
* bcd_in1=10000110 bcd_in2=10001000 cout=1 sum=01110100
* bcd_in1=10000110 bcd_in2=10001001 cout=1 sum=01110101
* bcd_in1=10000110 bcd_in2=10010000 cout=1 sum=01110110
* bcd_in1=10000110 bcd_in2=10010001 cout=1 sum=01110111
* bcd_in1=10000110 bcd_in2=10010010 cout=1 sum=01111000
* bcd_in1=10000110 bcd_in2=10010011 cout=1 sum=01111001
* bcd_in1=10000110 bcd_in2=10010100 cout=1 sum=10000000
* bcd_in1=10000110 bcd_in2=10010101 cout=1 sum=10000001
* bcd_in1=10000110 bcd_in2=10010110 cout=1 sum=10000010
* bcd_in1=10000110 bcd_in2=10010111 cout=1 sum=10000011
* bcd_in1=10000110 bcd_in2=10011000 cout=1 sum=10000100
* bcd_in1=10000110 bcd_in2=10011001 cout=1 sum=10000101
* bcd_in1=10000111 bcd_in2=00000000 cout=0 sum=10000111
* bcd_in1=10000111 bcd_in2=00000001 cout=0 sum=10001000
* bcd_in1=10000111 bcd_in2=00000010 cout=0 sum=10001001
* bcd_in1=10000111 bcd_in2=00000011 cout=0 sum=10010000
* bcd_in1=10000111 bcd_in2=00000100 cout=0 sum=10010001
* bcd_in1=10000111 bcd_in2=00000101 cout=0 sum=10010010
* bcd_in1=10000111 bcd_in2=00000110 cout=0 sum=10010011
* bcd_in1=10000111 bcd_in2=00000111 cout=0 sum=10010100
* bcd_in1=10000111 bcd_in2=00001000 cout=0 sum=10010101
* bcd_in1=10000111 bcd_in2=00001001 cout=0 sum=10010110
* bcd_in1=10000111 bcd_in2=00010000 cout=0 sum=10010111
* bcd_in1=10000111 bcd_in2=00010001 cout=0 sum=10011000
* bcd_in1=10000111 bcd_in2=00010010 cout=0 sum=10011001
* bcd_in1=10000111 bcd_in2=00010011 cout=1 sum=00000000
* bcd_in1=10000111 bcd_in2=00010100 cout=1 sum=00000001
* bcd_in1=10000111 bcd_in2=00010101 cout=1 sum=00000010
* bcd_in1=10000111 bcd_in2=00010110 cout=1 sum=00000011
* bcd_in1=10000111 bcd_in2=00010111 cout=1 sum=00000100
* bcd_in1=10000111 bcd_in2=00011000 cout=1 sum=00000101
* bcd_in1=10000111 bcd_in2=00011001 cout=1 sum=00000110
* bcd_in1=10000111 bcd_in2=00100000 cout=1 sum=00000111
* bcd_in1=10000111 bcd_in2=00100001 cout=1 sum=00001000
* bcd_in1=10000111 bcd_in2=00100010 cout=1 sum=00001001
* bcd_in1=10000111 bcd_in2=00100011 cout=1 sum=00010000
* bcd_in1=10000111 bcd_in2=00100100 cout=1 sum=00010001
* bcd_in1=10000111 bcd_in2=00100101 cout=1 sum=00010010
* bcd_in1=10000111 bcd_in2=00100110 cout=1 sum=00010011
* bcd_in1=10000111 bcd_in2=00100111 cout=1 sum=00010100
* bcd_in1=10000111 bcd_in2=00101000 cout=1 sum=00010101
* bcd_in1=10000111 bcd_in2=00101001 cout=1 sum=00010110
* bcd_in1=10000111 bcd_in2=00110000 cout=1 sum=00010111
* bcd_in1=10000111 bcd_in2=00110001 cout=1 sum=00011000
* bcd_in1=10000111 bcd_in2=00110010 cout=1 sum=00011001
* bcd_in1=10000111 bcd_in2=00110011 cout=1 sum=00100000
* bcd_in1=10000111 bcd_in2=00110100 cout=1 sum=00100001
* bcd_in1=10000111 bcd_in2=00110101 cout=1 sum=00100010
* bcd_in1=10000111 bcd_in2=00110110 cout=1 sum=00100011
* bcd_in1=10000111 bcd_in2=00110111 cout=1 sum=00100100
* bcd_in1=10000111 bcd_in2=00111000 cout=1 sum=00100101
* bcd_in1=10000111 bcd_in2=00111001 cout=1 sum=00100110
* bcd_in1=10000111 bcd_in2=01000000 cout=1 sum=00100111
* bcd_in1=10000111 bcd_in2=01000001 cout=1 sum=00101000
* bcd_in1=10000111 bcd_in2=01000010 cout=1 sum=00101001
* bcd_in1=10000111 bcd_in2=01000011 cout=1 sum=00110000
* bcd_in1=10000111 bcd_in2=01000100 cout=1 sum=00110001
* bcd_in1=10000111 bcd_in2=01000101 cout=1 sum=00110010
* bcd_in1=10000111 bcd_in2=01000110 cout=1 sum=00110011
* bcd_in1=10000111 bcd_in2=01000111 cout=1 sum=00110100
* bcd_in1=10000111 bcd_in2=01001000 cout=1 sum=00110101
* bcd_in1=10000111 bcd_in2=01001001 cout=1 sum=00110110
* bcd_in1=10000111 bcd_in2=01010000 cout=1 sum=00110111
* bcd_in1=10000111 bcd_in2=01010001 cout=1 sum=00111000
* bcd_in1=10000111 bcd_in2=01010010 cout=1 sum=00111001
* bcd_in1=10000111 bcd_in2=01010011 cout=1 sum=01000000
* bcd_in1=10000111 bcd_in2=01010100 cout=1 sum=01000001
* bcd_in1=10000111 bcd_in2=01010101 cout=1 sum=01000010
* bcd_in1=10000111 bcd_in2=01010110 cout=1 sum=01000011
* bcd_in1=10000111 bcd_in2=01010111 cout=1 sum=01000100
* bcd_in1=10000111 bcd_in2=01011000 cout=1 sum=01000101
* bcd_in1=10000111 bcd_in2=01011001 cout=1 sum=01000110
* bcd_in1=10000111 bcd_in2=01100000 cout=1 sum=01000111
* bcd_in1=10000111 bcd_in2=01100001 cout=1 sum=01001000
* bcd_in1=10000111 bcd_in2=01100010 cout=1 sum=01001001
* bcd_in1=10000111 bcd_in2=01100011 cout=1 sum=01010000
* bcd_in1=10000111 bcd_in2=01100100 cout=1 sum=01010001
* bcd_in1=10000111 bcd_in2=01100101 cout=1 sum=01010010
* bcd_in1=10000111 bcd_in2=01100110 cout=1 sum=01010011
* bcd_in1=10000111 bcd_in2=01100111 cout=1 sum=01010100
* bcd_in1=10000111 bcd_in2=01101000 cout=1 sum=01010101
* bcd_in1=10000111 bcd_in2=01101001 cout=1 sum=01010110
* bcd_in1=10000111 bcd_in2=01110000 cout=1 sum=01010111
* bcd_in1=10000111 bcd_in2=01110001 cout=1 sum=01011000
* bcd_in1=10000111 bcd_in2=01110010 cout=1 sum=01011001
* bcd_in1=10000111 bcd_in2=01110011 cout=1 sum=01100000
* bcd_in1=10000111 bcd_in2=01110100 cout=1 sum=01100001
* bcd_in1=10000111 bcd_in2=01110101 cout=1 sum=01100010
* bcd_in1=10000111 bcd_in2=01110110 cout=1 sum=01100011
* bcd_in1=10000111 bcd_in2=01110111 cout=1 sum=01100100
* bcd_in1=10000111 bcd_in2=01111000 cout=1 sum=01100101
* bcd_in1=10000111 bcd_in2=01111001 cout=1 sum=01100110
* bcd_in1=10000111 bcd_in2=10000000 cout=1 sum=01100111
* bcd_in1=10000111 bcd_in2=10000001 cout=1 sum=01101000
* bcd_in1=10000111 bcd_in2=10000010 cout=1 sum=01101001
* bcd_in1=10000111 bcd_in2=10000011 cout=1 sum=01110000
* bcd_in1=10000111 bcd_in2=10000100 cout=1 sum=01110001
* bcd_in1=10000111 bcd_in2=10000101 cout=1 sum=01110010
* bcd_in1=10000111 bcd_in2=10000110 cout=1 sum=01110011
* bcd_in1=10000111 bcd_in2=10000111 cout=1 sum=01110100
* bcd_in1=10000111 bcd_in2=10001000 cout=1 sum=01110101
* bcd_in1=10000111 bcd_in2=10001001 cout=1 sum=01110110
* bcd_in1=10000111 bcd_in2=10010000 cout=1 sum=01110111
* bcd_in1=10000111 bcd_in2=10010001 cout=1 sum=01111000
* bcd_in1=10000111 bcd_in2=10010010 cout=1 sum=01111001
* bcd_in1=10000111 bcd_in2=10010011 cout=1 sum=10000000
* bcd_in1=10000111 bcd_in2=10010100 cout=1 sum=10000001
* bcd_in1=10000111 bcd_in2=10010101 cout=1 sum=10000010
* bcd_in1=10000111 bcd_in2=10010110 cout=1 sum=10000011
* bcd_in1=10000111 bcd_in2=10010111 cout=1 sum=10000100
* bcd_in1=10000111 bcd_in2=10011000 cout=1 sum=10000101
* bcd_in1=10000111 bcd_in2=10011001 cout=1 sum=10000110
* bcd_in1=10001000 bcd_in2=00000000 cout=0 sum=10001000
* bcd_in1=10001000 bcd_in2=00000001 cout=0 sum=10001001
* bcd_in1=10001000 bcd_in2=00000010 cout=0 sum=10010000
* bcd_in1=10001000 bcd_in2=00000011 cout=0 sum=10010001
* bcd_in1=10001000 bcd_in2=00000100 cout=0 sum=10010010
* bcd_in1=10001000 bcd_in2=00000101 cout=0 sum=10010011
* bcd_in1=10001000 bcd_in2=00000110 cout=0 sum=10010100
* bcd_in1=10001000 bcd_in2=00000111 cout=0 sum=10010101
* bcd_in1=10001000 bcd_in2=00001000 cout=0 sum=10010110
* bcd_in1=10001000 bcd_in2=00001001 cout=0 sum=10010111
* bcd_in1=10001000 bcd_in2=00010000 cout=0 sum=10011000
* bcd_in1=10001000 bcd_in2=00010001 cout=0 sum=10011001
* bcd_in1=10001000 bcd_in2=00010010 cout=1 sum=00000000
* bcd_in1=10001000 bcd_in2=00010011 cout=1 sum=00000001
* bcd_in1=10001000 bcd_in2=00010100 cout=1 sum=00000010
* bcd_in1=10001000 bcd_in2=00010101 cout=1 sum=00000011
* bcd_in1=10001000 bcd_in2=00010110 cout=1 sum=00000100
* bcd_in1=10001000 bcd_in2=00010111 cout=1 sum=00000101
* bcd_in1=10001000 bcd_in2=00011000 cout=1 sum=00000110
* bcd_in1=10001000 bcd_in2=00011001 cout=1 sum=00000111
* bcd_in1=10001000 bcd_in2=00100000 cout=1 sum=00001000
* bcd_in1=10001000 bcd_in2=00100001 cout=1 sum=00001001
* bcd_in1=10001000 bcd_in2=00100010 cout=1 sum=00010000
* bcd_in1=10001000 bcd_in2=00100011 cout=1 sum=00010001
* bcd_in1=10001000 bcd_in2=00100100 cout=1 sum=00010010
* bcd_in1=10001000 bcd_in2=00100101 cout=1 sum=00010011
* bcd_in1=10001000 bcd_in2=00100110 cout=1 sum=00010100
* bcd_in1=10001000 bcd_in2=00100111 cout=1 sum=00010101
* bcd_in1=10001000 bcd_in2=00101000 cout=1 sum=00010110
* bcd_in1=10001000 bcd_in2=00101001 cout=1 sum=00010111
* bcd_in1=10001000 bcd_in2=00110000 cout=1 sum=00011000
* bcd_in1=10001000 bcd_in2=00110001 cout=1 sum=00011001
* bcd_in1=10001000 bcd_in2=00110010 cout=1 sum=00100000
* bcd_in1=10001000 bcd_in2=00110011 cout=1 sum=00100001
* bcd_in1=10001000 bcd_in2=00110100 cout=1 sum=00100010
* bcd_in1=10001000 bcd_in2=00110101 cout=1 sum=00100011
* bcd_in1=10001000 bcd_in2=00110110 cout=1 sum=00100100
* bcd_in1=10001000 bcd_in2=00110111 cout=1 sum=00100101
* bcd_in1=10001000 bcd_in2=00111000 cout=1 sum=00100110
* bcd_in1=10001000 bcd_in2=00111001 cout=1 sum=00100111
* bcd_in1=10001000 bcd_in2=01000000 cout=1 sum=00101000
* bcd_in1=10001000 bcd_in2=01000001 cout=1 sum=00101001
* bcd_in1=10001000 bcd_in2=01000010 cout=1 sum=00110000
* bcd_in1=10001000 bcd_in2=01000011 cout=1 sum=00110001
* bcd_in1=10001000 bcd_in2=01000100 cout=1 sum=00110010
* bcd_in1=10001000 bcd_in2=01000101 cout=1 sum=00110011
* bcd_in1=10001000 bcd_in2=01000110 cout=1 sum=00110100
* bcd_in1=10001000 bcd_in2=01000111 cout=1 sum=00110101
* bcd_in1=10001000 bcd_in2=01001000 cout=1 sum=00110110
* bcd_in1=10001000 bcd_in2=01001001 cout=1 sum=00110111
* bcd_in1=10001000 bcd_in2=01010000 cout=1 sum=00111000
* bcd_in1=10001000 bcd_in2=01010001 cout=1 sum=00111001
* bcd_in1=10001000 bcd_in2=01010010 cout=1 sum=01000000
* bcd_in1=10001000 bcd_in2=01010011 cout=1 sum=01000001
* bcd_in1=10001000 bcd_in2=01010100 cout=1 sum=01000010
* bcd_in1=10001000 bcd_in2=01010101 cout=1 sum=01000011
* bcd_in1=10001000 bcd_in2=01010110 cout=1 sum=01000100
* bcd_in1=10001000 bcd_in2=01010111 cout=1 sum=01000101
* bcd_in1=10001000 bcd_in2=01011000 cout=1 sum=01000110
* bcd_in1=10001000 bcd_in2=01011001 cout=1 sum=01000111
* bcd_in1=10001000 bcd_in2=01100000 cout=1 sum=01001000
* bcd_in1=10001000 bcd_in2=01100001 cout=1 sum=01001001
* bcd_in1=10001000 bcd_in2=01100010 cout=1 sum=01010000
* bcd_in1=10001000 bcd_in2=01100011 cout=1 sum=01010001
* bcd_in1=10001000 bcd_in2=01100100 cout=1 sum=01010010
* bcd_in1=10001000 bcd_in2=01100101 cout=1 sum=01010011
* bcd_in1=10001000 bcd_in2=01100110 cout=1 sum=01010100
* bcd_in1=10001000 bcd_in2=01100111 cout=1 sum=01010101
* bcd_in1=10001000 bcd_in2=01101000 cout=1 sum=01010110
* bcd_in1=10001000 bcd_in2=01101001 cout=1 sum=01010111
* bcd_in1=10001000 bcd_in2=01110000 cout=1 sum=01011000
* bcd_in1=10001000 bcd_in2=01110001 cout=1 sum=01011001
* bcd_in1=10001000 bcd_in2=01110010 cout=1 sum=01100000
* bcd_in1=10001000 bcd_in2=01110011 cout=1 sum=01100001
* bcd_in1=10001000 bcd_in2=01110100 cout=1 sum=01100010
* bcd_in1=10001000 bcd_in2=01110101 cout=1 sum=01100011
* bcd_in1=10001000 bcd_in2=01110110 cout=1 sum=01100100
* bcd_in1=10001000 bcd_in2=01110111 cout=1 sum=01100101
* bcd_in1=10001000 bcd_in2=01111000 cout=1 sum=01100110
* bcd_in1=10001000 bcd_in2=01111001 cout=1 sum=01100111
* bcd_in1=10001000 bcd_in2=10000000 cout=1 sum=01101000
* bcd_in1=10001000 bcd_in2=10000001 cout=1 sum=01101001
* bcd_in1=10001000 bcd_in2=10000010 cout=1 sum=01110000
* bcd_in1=10001000 bcd_in2=10000011 cout=1 sum=01110001
* bcd_in1=10001000 bcd_in2=10000100 cout=1 sum=01110010
* bcd_in1=10001000 bcd_in2=10000101 cout=1 sum=01110011
* bcd_in1=10001000 bcd_in2=10000110 cout=1 sum=01110100
* bcd_in1=10001000 bcd_in2=10000111 cout=1 sum=01110101
* bcd_in1=10001000 bcd_in2=10001000 cout=1 sum=01110110
* bcd_in1=10001000 bcd_in2=10001001 cout=1 sum=01110111
* bcd_in1=10001000 bcd_in2=10010000 cout=1 sum=01111000
* bcd_in1=10001000 bcd_in2=10010001 cout=1 sum=01111001
* bcd_in1=10001000 bcd_in2=10010010 cout=1 sum=10000000
* bcd_in1=10001000 bcd_in2=10010011 cout=1 sum=10000001
* bcd_in1=10001000 bcd_in2=10010100 cout=1 sum=10000010
* bcd_in1=10001000 bcd_in2=10010101 cout=1 sum=10000011
* bcd_in1=10001000 bcd_in2=10010110 cout=1 sum=10000100
* bcd_in1=10001000 bcd_in2=10010111 cout=1 sum=10000101
* bcd_in1=10001000 bcd_in2=10011000 cout=1 sum=10000110
* bcd_in1=10001000 bcd_in2=10011001 cout=1 sum=10000111
* bcd_in1=10001001 bcd_in2=00000000 cout=0 sum=10001001
* bcd_in1=10001001 bcd_in2=00000001 cout=0 sum=10010000
* bcd_in1=10001001 bcd_in2=00000010 cout=0 sum=10010001
* bcd_in1=10001001 bcd_in2=00000011 cout=0 sum=10010010
* bcd_in1=10001001 bcd_in2=00000100 cout=0 sum=10010011
* bcd_in1=10001001 bcd_in2=00000101 cout=0 sum=10010100
* bcd_in1=10001001 bcd_in2=00000110 cout=0 sum=10010101
* bcd_in1=10001001 bcd_in2=00000111 cout=0 sum=10010110
* bcd_in1=10001001 bcd_in2=00001000 cout=0 sum=10010111
* bcd_in1=10001001 bcd_in2=00001001 cout=0 sum=10011000
* bcd_in1=10001001 bcd_in2=00010000 cout=0 sum=10011001
* bcd_in1=10001001 bcd_in2=00010001 cout=1 sum=00000000
* bcd_in1=10001001 bcd_in2=00010010 cout=1 sum=00000001
* bcd_in1=10001001 bcd_in2=00010011 cout=1 sum=00000010
* bcd_in1=10001001 bcd_in2=00010100 cout=1 sum=00000011
* bcd_in1=10001001 bcd_in2=00010101 cout=1 sum=00000100
* bcd_in1=10001001 bcd_in2=00010110 cout=1 sum=00000101
* bcd_in1=10001001 bcd_in2=00010111 cout=1 sum=00000110
* bcd_in1=10001001 bcd_in2=00011000 cout=1 sum=00000111
* bcd_in1=10001001 bcd_in2=00011001 cout=1 sum=00001000
* bcd_in1=10001001 bcd_in2=00100000 cout=1 sum=00001001
* bcd_in1=10001001 bcd_in2=00100001 cout=1 sum=00010000
* bcd_in1=10001001 bcd_in2=00100010 cout=1 sum=00010001
* bcd_in1=10001001 bcd_in2=00100011 cout=1 sum=00010010
* bcd_in1=10001001 bcd_in2=00100100 cout=1 sum=00010011
* bcd_in1=10001001 bcd_in2=00100101 cout=1 sum=00010100
* bcd_in1=10001001 bcd_in2=00100110 cout=1 sum=00010101
* bcd_in1=10001001 bcd_in2=00100111 cout=1 sum=00010110
* bcd_in1=10001001 bcd_in2=00101000 cout=1 sum=00010111
* bcd_in1=10001001 bcd_in2=00101001 cout=1 sum=00011000
* bcd_in1=10001001 bcd_in2=00110000 cout=1 sum=00011001
* bcd_in1=10001001 bcd_in2=00110001 cout=1 sum=00100000
* bcd_in1=10001001 bcd_in2=00110010 cout=1 sum=00100001
* bcd_in1=10001001 bcd_in2=00110011 cout=1 sum=00100010
* bcd_in1=10001001 bcd_in2=00110100 cout=1 sum=00100011
* bcd_in1=10001001 bcd_in2=00110101 cout=1 sum=00100100
* bcd_in1=10001001 bcd_in2=00110110 cout=1 sum=00100101
* bcd_in1=10001001 bcd_in2=00110111 cout=1 sum=00100110
* bcd_in1=10001001 bcd_in2=00111000 cout=1 sum=00100111
* bcd_in1=10001001 bcd_in2=00111001 cout=1 sum=00101000
* bcd_in1=10001001 bcd_in2=01000000 cout=1 sum=00101001
* bcd_in1=10001001 bcd_in2=01000001 cout=1 sum=00110000
* bcd_in1=10001001 bcd_in2=01000010 cout=1 sum=00110001
* bcd_in1=10001001 bcd_in2=01000011 cout=1 sum=00110010
* bcd_in1=10001001 bcd_in2=01000100 cout=1 sum=00110011
* bcd_in1=10001001 bcd_in2=01000101 cout=1 sum=00110100
* bcd_in1=10001001 bcd_in2=01000110 cout=1 sum=00110101
* bcd_in1=10001001 bcd_in2=01000111 cout=1 sum=00110110
* bcd_in1=10001001 bcd_in2=01001000 cout=1 sum=00110111
* bcd_in1=10001001 bcd_in2=01001001 cout=1 sum=00111000
* bcd_in1=10001001 bcd_in2=01010000 cout=1 sum=00111001
* bcd_in1=10001001 bcd_in2=01010001 cout=1 sum=01000000
* bcd_in1=10001001 bcd_in2=01010010 cout=1 sum=01000001
* bcd_in1=10001001 bcd_in2=01010011 cout=1 sum=01000010
* bcd_in1=10001001 bcd_in2=01010100 cout=1 sum=01000011
* bcd_in1=10001001 bcd_in2=01010101 cout=1 sum=01000100
* bcd_in1=10001001 bcd_in2=01010110 cout=1 sum=01000101
* bcd_in1=10001001 bcd_in2=01010111 cout=1 sum=01000110
* bcd_in1=10001001 bcd_in2=01011000 cout=1 sum=01000111
* bcd_in1=10001001 bcd_in2=01011001 cout=1 sum=01001000
* bcd_in1=10001001 bcd_in2=01100000 cout=1 sum=01001001
* bcd_in1=10001001 bcd_in2=01100001 cout=1 sum=01010000
* bcd_in1=10001001 bcd_in2=01100010 cout=1 sum=01010001
* bcd_in1=10001001 bcd_in2=01100011 cout=1 sum=01010010
* bcd_in1=10001001 bcd_in2=01100100 cout=1 sum=01010011
* bcd_in1=10001001 bcd_in2=01100101 cout=1 sum=01010100
* bcd_in1=10001001 bcd_in2=01100110 cout=1 sum=01010101
* bcd_in1=10001001 bcd_in2=01100111 cout=1 sum=01010110
* bcd_in1=10001001 bcd_in2=01101000 cout=1 sum=01010111
* bcd_in1=10001001 bcd_in2=01101001 cout=1 sum=01011000
* bcd_in1=10001001 bcd_in2=01110000 cout=1 sum=01011001
* bcd_in1=10001001 bcd_in2=01110001 cout=1 sum=01100000
* bcd_in1=10001001 bcd_in2=01110010 cout=1 sum=01100001
* bcd_in1=10001001 bcd_in2=01110011 cout=1 sum=01100010
* bcd_in1=10001001 bcd_in2=01110100 cout=1 sum=01100011
* bcd_in1=10001001 bcd_in2=01110101 cout=1 sum=01100100
* bcd_in1=10001001 bcd_in2=01110110 cout=1 sum=01100101
* bcd_in1=10001001 bcd_in2=01110111 cout=1 sum=01100110
* bcd_in1=10001001 bcd_in2=01111000 cout=1 sum=01100111
* bcd_in1=10001001 bcd_in2=01111001 cout=1 sum=01101000
* bcd_in1=10001001 bcd_in2=10000000 cout=1 sum=01101001
* bcd_in1=10001001 bcd_in2=10000001 cout=1 sum=01110000
* bcd_in1=10001001 bcd_in2=10000010 cout=1 sum=01110001
* bcd_in1=10001001 bcd_in2=10000011 cout=1 sum=01110010
* bcd_in1=10001001 bcd_in2=10000100 cout=1 sum=01110011
* bcd_in1=10001001 bcd_in2=10000101 cout=1 sum=01110100
* bcd_in1=10001001 bcd_in2=10000110 cout=1 sum=01110101
* bcd_in1=10001001 bcd_in2=10000111 cout=1 sum=01110110
* bcd_in1=10001001 bcd_in2=10001000 cout=1 sum=01110111
* bcd_in1=10001001 bcd_in2=10001001 cout=1 sum=01111000
* bcd_in1=10001001 bcd_in2=10010000 cout=1 sum=01111001
* bcd_in1=10001001 bcd_in2=10010001 cout=1 sum=10000000
* bcd_in1=10001001 bcd_in2=10010010 cout=1 sum=10000001
* bcd_in1=10001001 bcd_in2=10010011 cout=1 sum=10000010
* bcd_in1=10001001 bcd_in2=10010100 cout=1 sum=10000011
* bcd_in1=10001001 bcd_in2=10010101 cout=1 sum=10000100
* bcd_in1=10001001 bcd_in2=10010110 cout=1 sum=10000101
* bcd_in1=10001001 bcd_in2=10010111 cout=1 sum=10000110
* bcd_in1=10001001 bcd_in2=10011000 cout=1 sum=10000111
* bcd_in1=10001001 bcd_in2=10011001 cout=1 sum=10001000
* bcd_in1=10010000 bcd_in2=00000000 cout=0 sum=10010000
* bcd_in1=10010000 bcd_in2=00000001 cout=0 sum=10010001
* bcd_in1=10010000 bcd_in2=00000010 cout=0 sum=10010010
* bcd_in1=10010000 bcd_in2=00000011 cout=0 sum=10010011
* bcd_in1=10010000 bcd_in2=00000100 cout=0 sum=10010100
* bcd_in1=10010000 bcd_in2=00000101 cout=0 sum=10010101
* bcd_in1=10010000 bcd_in2=00000110 cout=0 sum=10010110
* bcd_in1=10010000 bcd_in2=00000111 cout=0 sum=10010111
* bcd_in1=10010000 bcd_in2=00001000 cout=0 sum=10011000
* bcd_in1=10010000 bcd_in2=00001001 cout=0 sum=10011001
* bcd_in1=10010000 bcd_in2=00010000 cout=1 sum=00000000
* bcd_in1=10010000 bcd_in2=00010001 cout=1 sum=00000001
* bcd_in1=10010000 bcd_in2=00010010 cout=1 sum=00000010
* bcd_in1=10010000 bcd_in2=00010011 cout=1 sum=00000011
* bcd_in1=10010000 bcd_in2=00010100 cout=1 sum=00000100
* bcd_in1=10010000 bcd_in2=00010101 cout=1 sum=00000101
* bcd_in1=10010000 bcd_in2=00010110 cout=1 sum=00000110
* bcd_in1=10010000 bcd_in2=00010111 cout=1 sum=00000111
* bcd_in1=10010000 bcd_in2=00011000 cout=1 sum=00001000
* bcd_in1=10010000 bcd_in2=00011001 cout=1 sum=00001001
* bcd_in1=10010000 bcd_in2=00100000 cout=1 sum=00010000
* bcd_in1=10010000 bcd_in2=00100001 cout=1 sum=00010001
* bcd_in1=10010000 bcd_in2=00100010 cout=1 sum=00010010
* bcd_in1=10010000 bcd_in2=00100011 cout=1 sum=00010011
* bcd_in1=10010000 bcd_in2=00100100 cout=1 sum=00010100
* bcd_in1=10010000 bcd_in2=00100101 cout=1 sum=00010101
* bcd_in1=10010000 bcd_in2=00100110 cout=1 sum=00010110
* bcd_in1=10010000 bcd_in2=00100111 cout=1 sum=00010111
* bcd_in1=10010000 bcd_in2=00101000 cout=1 sum=00011000
* bcd_in1=10010000 bcd_in2=00101001 cout=1 sum=00011001
* bcd_in1=10010000 bcd_in2=00110000 cout=1 sum=00100000
* bcd_in1=10010000 bcd_in2=00110001 cout=1 sum=00100001
* bcd_in1=10010000 bcd_in2=00110010 cout=1 sum=00100010
* bcd_in1=10010000 bcd_in2=00110011 cout=1 sum=00100011
* bcd_in1=10010000 bcd_in2=00110100 cout=1 sum=00100100
* bcd_in1=10010000 bcd_in2=00110101 cout=1 sum=00100101
* bcd_in1=10010000 bcd_in2=00110110 cout=1 sum=00100110
* bcd_in1=10010000 bcd_in2=00110111 cout=1 sum=00100111
* bcd_in1=10010000 bcd_in2=00111000 cout=1 sum=00101000
* bcd_in1=10010000 bcd_in2=00111001 cout=1 sum=00101001
* bcd_in1=10010000 bcd_in2=01000000 cout=1 sum=00110000
* bcd_in1=10010000 bcd_in2=01000001 cout=1 sum=00110001
* bcd_in1=10010000 bcd_in2=01000010 cout=1 sum=00110010
* bcd_in1=10010000 bcd_in2=01000011 cout=1 sum=00110011
* bcd_in1=10010000 bcd_in2=01000100 cout=1 sum=00110100
* bcd_in1=10010000 bcd_in2=01000101 cout=1 sum=00110101
* bcd_in1=10010000 bcd_in2=01000110 cout=1 sum=00110110
* bcd_in1=10010000 bcd_in2=01000111 cout=1 sum=00110111
* bcd_in1=10010000 bcd_in2=01001000 cout=1 sum=00111000
* bcd_in1=10010000 bcd_in2=01001001 cout=1 sum=00111001
* bcd_in1=10010000 bcd_in2=01010000 cout=1 sum=01000000
* bcd_in1=10010000 bcd_in2=01010001 cout=1 sum=01000001
* bcd_in1=10010000 bcd_in2=01010010 cout=1 sum=01000010
* bcd_in1=10010000 bcd_in2=01010011 cout=1 sum=01000011
* bcd_in1=10010000 bcd_in2=01010100 cout=1 sum=01000100
* bcd_in1=10010000 bcd_in2=01010101 cout=1 sum=01000101
* bcd_in1=10010000 bcd_in2=01010110 cout=1 sum=01000110
* bcd_in1=10010000 bcd_in2=01010111 cout=1 sum=01000111
* bcd_in1=10010000 bcd_in2=01011000 cout=1 sum=01001000
* bcd_in1=10010000 bcd_in2=01011001 cout=1 sum=01001001
* bcd_in1=10010000 bcd_in2=01100000 cout=1 sum=01010000
* bcd_in1=10010000 bcd_in2=01100001 cout=1 sum=01010001
* bcd_in1=10010000 bcd_in2=01100010 cout=1 sum=01010010
* bcd_in1=10010000 bcd_in2=01100011 cout=1 sum=01010011
* bcd_in1=10010000 bcd_in2=01100100 cout=1 sum=01010100
* bcd_in1=10010000 bcd_in2=01100101 cout=1 sum=01010101
* bcd_in1=10010000 bcd_in2=01100110 cout=1 sum=01010110
* bcd_in1=10010000 bcd_in2=01100111 cout=1 sum=01010111
* bcd_in1=10010000 bcd_in2=01101000 cout=1 sum=01011000
* bcd_in1=10010000 bcd_in2=01101001 cout=1 sum=01011001
* bcd_in1=10010000 bcd_in2=01110000 cout=1 sum=01100000
* bcd_in1=10010000 bcd_in2=01110001 cout=1 sum=01100001
* bcd_in1=10010000 bcd_in2=01110010 cout=1 sum=01100010
* bcd_in1=10010000 bcd_in2=01110011 cout=1 sum=01100011
* bcd_in1=10010000 bcd_in2=01110100 cout=1 sum=01100100
* bcd_in1=10010000 bcd_in2=01110101 cout=1 sum=01100101
* bcd_in1=10010000 bcd_in2=01110110 cout=1 sum=01100110
* bcd_in1=10010000 bcd_in2=01110111 cout=1 sum=01100111
* bcd_in1=10010000 bcd_in2=01111000 cout=1 sum=01101000
* bcd_in1=10010000 bcd_in2=01111001 cout=1 sum=01101001
* bcd_in1=10010000 bcd_in2=10000000 cout=1 sum=01110000
* bcd_in1=10010000 bcd_in2=10000001 cout=1 sum=01110001
* bcd_in1=10010000 bcd_in2=10000010 cout=1 sum=01110010
* bcd_in1=10010000 bcd_in2=10000011 cout=1 sum=01110011
* bcd_in1=10010000 bcd_in2=10000100 cout=1 sum=01110100
* bcd_in1=10010000 bcd_in2=10000101 cout=1 sum=01110101
* bcd_in1=10010000 bcd_in2=10000110 cout=1 sum=01110110
* bcd_in1=10010000 bcd_in2=10000111 cout=1 sum=01110111
* bcd_in1=10010000 bcd_in2=10001000 cout=1 sum=01111000
* bcd_in1=10010000 bcd_in2=10001001 cout=1 sum=01111001
* bcd_in1=10010000 bcd_in2=10010000 cout=1 sum=10000000
* bcd_in1=10010000 bcd_in2=10010001 cout=1 sum=10000001
* bcd_in1=10010000 bcd_in2=10010010 cout=1 sum=10000010
* bcd_in1=10010000 bcd_in2=10010011 cout=1 sum=10000011
* bcd_in1=10010000 bcd_in2=10010100 cout=1 sum=10000100
* bcd_in1=10010000 bcd_in2=10010101 cout=1 sum=10000101
* bcd_in1=10010000 bcd_in2=10010110 cout=1 sum=10000110
* bcd_in1=10010000 bcd_in2=10010111 cout=1 sum=10000111
* bcd_in1=10010000 bcd_in2=10011000 cout=1 sum=10001000
* bcd_in1=10010000 bcd_in2=10011001 cout=1 sum=10001001
* bcd_in1=10010001 bcd_in2=00000000 cout=0 sum=10010001
* bcd_in1=10010001 bcd_in2=00000001 cout=0 sum=10010010
* bcd_in1=10010001 bcd_in2=00000010 cout=0 sum=10010011
* bcd_in1=10010001 bcd_in2=00000011 cout=0 sum=10010100
* bcd_in1=10010001 bcd_in2=00000100 cout=0 sum=10010101
* bcd_in1=10010001 bcd_in2=00000101 cout=0 sum=10010110
* bcd_in1=10010001 bcd_in2=00000110 cout=0 sum=10010111
* bcd_in1=10010001 bcd_in2=00000111 cout=0 sum=10011000
* bcd_in1=10010001 bcd_in2=00001000 cout=0 sum=10011001
* bcd_in1=10010001 bcd_in2=00001001 cout=1 sum=00000000
* bcd_in1=10010001 bcd_in2=00010000 cout=1 sum=00000001
* bcd_in1=10010001 bcd_in2=00010001 cout=1 sum=00000010
* bcd_in1=10010001 bcd_in2=00010010 cout=1 sum=00000011
* bcd_in1=10010001 bcd_in2=00010011 cout=1 sum=00000100
* bcd_in1=10010001 bcd_in2=00010100 cout=1 sum=00000101
* bcd_in1=10010001 bcd_in2=00010101 cout=1 sum=00000110
* bcd_in1=10010001 bcd_in2=00010110 cout=1 sum=00000111
* bcd_in1=10010001 bcd_in2=00010111 cout=1 sum=00001000
* bcd_in1=10010001 bcd_in2=00011000 cout=1 sum=00001001
* bcd_in1=10010001 bcd_in2=00011001 cout=1 sum=00010000
* bcd_in1=10010001 bcd_in2=00100000 cout=1 sum=00010001
* bcd_in1=10010001 bcd_in2=00100001 cout=1 sum=00010010
* bcd_in1=10010001 bcd_in2=00100010 cout=1 sum=00010011
* bcd_in1=10010001 bcd_in2=00100011 cout=1 sum=00010100
* bcd_in1=10010001 bcd_in2=00100100 cout=1 sum=00010101
* bcd_in1=10010001 bcd_in2=00100101 cout=1 sum=00010110
* bcd_in1=10010001 bcd_in2=00100110 cout=1 sum=00010111
* bcd_in1=10010001 bcd_in2=00100111 cout=1 sum=00011000
* bcd_in1=10010001 bcd_in2=00101000 cout=1 sum=00011001
* bcd_in1=10010001 bcd_in2=00101001 cout=1 sum=00100000
* bcd_in1=10010001 bcd_in2=00110000 cout=1 sum=00100001
* bcd_in1=10010001 bcd_in2=00110001 cout=1 sum=00100010
* bcd_in1=10010001 bcd_in2=00110010 cout=1 sum=00100011
* bcd_in1=10010001 bcd_in2=00110011 cout=1 sum=00100100
* bcd_in1=10010001 bcd_in2=00110100 cout=1 sum=00100101
* bcd_in1=10010001 bcd_in2=00110101 cout=1 sum=00100110
* bcd_in1=10010001 bcd_in2=00110110 cout=1 sum=00100111
* bcd_in1=10010001 bcd_in2=00110111 cout=1 sum=00101000
* bcd_in1=10010001 bcd_in2=00111000 cout=1 sum=00101001
* bcd_in1=10010001 bcd_in2=00111001 cout=1 sum=00110000
* bcd_in1=10010001 bcd_in2=01000000 cout=1 sum=00110001
* bcd_in1=10010001 bcd_in2=01000001 cout=1 sum=00110010
* bcd_in1=10010001 bcd_in2=01000010 cout=1 sum=00110011
* bcd_in1=10010001 bcd_in2=01000011 cout=1 sum=00110100
* bcd_in1=10010001 bcd_in2=01000100 cout=1 sum=00110101
* bcd_in1=10010001 bcd_in2=01000101 cout=1 sum=00110110
* bcd_in1=10010001 bcd_in2=01000110 cout=1 sum=00110111
* bcd_in1=10010001 bcd_in2=01000111 cout=1 sum=00111000
* bcd_in1=10010001 bcd_in2=01001000 cout=1 sum=00111001
* bcd_in1=10010001 bcd_in2=01001001 cout=1 sum=01000000
* bcd_in1=10010001 bcd_in2=01010000 cout=1 sum=01000001
* bcd_in1=10010001 bcd_in2=01010001 cout=1 sum=01000010
* bcd_in1=10010001 bcd_in2=01010010 cout=1 sum=01000011
* bcd_in1=10010001 bcd_in2=01010011 cout=1 sum=01000100
* bcd_in1=10010001 bcd_in2=01010100 cout=1 sum=01000101
* bcd_in1=10010001 bcd_in2=01010101 cout=1 sum=01000110
* bcd_in1=10010001 bcd_in2=01010110 cout=1 sum=01000111
* bcd_in1=10010001 bcd_in2=01010111 cout=1 sum=01001000
* bcd_in1=10010001 bcd_in2=01011000 cout=1 sum=01001001
* bcd_in1=10010001 bcd_in2=01011001 cout=1 sum=01010000
* bcd_in1=10010001 bcd_in2=01100000 cout=1 sum=01010001
* bcd_in1=10010001 bcd_in2=01100001 cout=1 sum=01010010
* bcd_in1=10010001 bcd_in2=01100010 cout=1 sum=01010011
* bcd_in1=10010001 bcd_in2=01100011 cout=1 sum=01010100
* bcd_in1=10010001 bcd_in2=01100100 cout=1 sum=01010101
* bcd_in1=10010001 bcd_in2=01100101 cout=1 sum=01010110
* bcd_in1=10010001 bcd_in2=01100110 cout=1 sum=01010111
* bcd_in1=10010001 bcd_in2=01100111 cout=1 sum=01011000
* bcd_in1=10010001 bcd_in2=01101000 cout=1 sum=01011001
* bcd_in1=10010001 bcd_in2=01101001 cout=1 sum=01100000
* bcd_in1=10010001 bcd_in2=01110000 cout=1 sum=01100001
* bcd_in1=10010001 bcd_in2=01110001 cout=1 sum=01100010
* bcd_in1=10010001 bcd_in2=01110010 cout=1 sum=01100011
* bcd_in1=10010001 bcd_in2=01110011 cout=1 sum=01100100
* bcd_in1=10010001 bcd_in2=01110100 cout=1 sum=01100101
* bcd_in1=10010001 bcd_in2=01110101 cout=1 sum=01100110
* bcd_in1=10010001 bcd_in2=01110110 cout=1 sum=01100111
* bcd_in1=10010001 bcd_in2=01110111 cout=1 sum=01101000
* bcd_in1=10010001 bcd_in2=01111000 cout=1 sum=01101001
* bcd_in1=10010001 bcd_in2=01111001 cout=1 sum=01110000
* bcd_in1=10010001 bcd_in2=10000000 cout=1 sum=01110001
* bcd_in1=10010001 bcd_in2=10000001 cout=1 sum=01110010
* bcd_in1=10010001 bcd_in2=10000010 cout=1 sum=01110011
* bcd_in1=10010001 bcd_in2=10000011 cout=1 sum=01110100
* bcd_in1=10010001 bcd_in2=10000100 cout=1 sum=01110101
* bcd_in1=10010001 bcd_in2=10000101 cout=1 sum=01110110
* bcd_in1=10010001 bcd_in2=10000110 cout=1 sum=01110111
* bcd_in1=10010001 bcd_in2=10000111 cout=1 sum=01111000
* bcd_in1=10010001 bcd_in2=10001000 cout=1 sum=01111001
* bcd_in1=10010001 bcd_in2=10001001 cout=1 sum=10000000
* bcd_in1=10010001 bcd_in2=10010000 cout=1 sum=10000001
* bcd_in1=10010001 bcd_in2=10010001 cout=1 sum=10000010
* bcd_in1=10010001 bcd_in2=10010010 cout=1 sum=10000011
* bcd_in1=10010001 bcd_in2=10010011 cout=1 sum=10000100
* bcd_in1=10010001 bcd_in2=10010100 cout=1 sum=10000101
* bcd_in1=10010001 bcd_in2=10010101 cout=1 sum=10000110
* bcd_in1=10010001 bcd_in2=10010110 cout=1 sum=10000111
* bcd_in1=10010001 bcd_in2=10010111 cout=1 sum=10001000
* bcd_in1=10010001 bcd_in2=10011000 cout=1 sum=10001001
* bcd_in1=10010001 bcd_in2=10011001 cout=1 sum=10010000
* bcd_in1=10010010 bcd_in2=00000000 cout=0 sum=10010010
* bcd_in1=10010010 bcd_in2=00000001 cout=0 sum=10010011
* bcd_in1=10010010 bcd_in2=00000010 cout=0 sum=10010100
* bcd_in1=10010010 bcd_in2=00000011 cout=0 sum=10010101
* bcd_in1=10010010 bcd_in2=00000100 cout=0 sum=10010110
* bcd_in1=10010010 bcd_in2=00000101 cout=0 sum=10010111
* bcd_in1=10010010 bcd_in2=00000110 cout=0 sum=10011000
* bcd_in1=10010010 bcd_in2=00000111 cout=0 sum=10011001
* bcd_in1=10010010 bcd_in2=00001000 cout=1 sum=00000000
* bcd_in1=10010010 bcd_in2=00001001 cout=1 sum=00000001
* bcd_in1=10010010 bcd_in2=00010000 cout=1 sum=00000010
* bcd_in1=10010010 bcd_in2=00010001 cout=1 sum=00000011
* bcd_in1=10010010 bcd_in2=00010010 cout=1 sum=00000100
* bcd_in1=10010010 bcd_in2=00010011 cout=1 sum=00000101
* bcd_in1=10010010 bcd_in2=00010100 cout=1 sum=00000110
* bcd_in1=10010010 bcd_in2=00010101 cout=1 sum=00000111
* bcd_in1=10010010 bcd_in2=00010110 cout=1 sum=00001000
* bcd_in1=10010010 bcd_in2=00010111 cout=1 sum=00001001
* bcd_in1=10010010 bcd_in2=00011000 cout=1 sum=00010000
* bcd_in1=10010010 bcd_in2=00011001 cout=1 sum=00010001
* bcd_in1=10010010 bcd_in2=00100000 cout=1 sum=00010010
* bcd_in1=10010010 bcd_in2=00100001 cout=1 sum=00010011
* bcd_in1=10010010 bcd_in2=00100010 cout=1 sum=00010100
* bcd_in1=10010010 bcd_in2=00100011 cout=1 sum=00010101
* bcd_in1=10010010 bcd_in2=00100100 cout=1 sum=00010110
* bcd_in1=10010010 bcd_in2=00100101 cout=1 sum=00010111
* bcd_in1=10010010 bcd_in2=00100110 cout=1 sum=00011000
* bcd_in1=10010010 bcd_in2=00100111 cout=1 sum=00011001
* bcd_in1=10010010 bcd_in2=00101000 cout=1 sum=00100000
* bcd_in1=10010010 bcd_in2=00101001 cout=1 sum=00100001
* bcd_in1=10010010 bcd_in2=00110000 cout=1 sum=00100010
* bcd_in1=10010010 bcd_in2=00110001 cout=1 sum=00100011
* bcd_in1=10010010 bcd_in2=00110010 cout=1 sum=00100100
* bcd_in1=10010010 bcd_in2=00110011 cout=1 sum=00100101
* bcd_in1=10010010 bcd_in2=00110100 cout=1 sum=00100110
* bcd_in1=10010010 bcd_in2=00110101 cout=1 sum=00100111
* bcd_in1=10010010 bcd_in2=00110110 cout=1 sum=00101000
* bcd_in1=10010010 bcd_in2=00110111 cout=1 sum=00101001
* bcd_in1=10010010 bcd_in2=00111000 cout=1 sum=00110000
* bcd_in1=10010010 bcd_in2=00111001 cout=1 sum=00110001
* bcd_in1=10010010 bcd_in2=01000000 cout=1 sum=00110010
* bcd_in1=10010010 bcd_in2=01000001 cout=1 sum=00110011
* bcd_in1=10010010 bcd_in2=01000010 cout=1 sum=00110100
* bcd_in1=10010010 bcd_in2=01000011 cout=1 sum=00110101
* bcd_in1=10010010 bcd_in2=01000100 cout=1 sum=00110110
* bcd_in1=10010010 bcd_in2=01000101 cout=1 sum=00110111
* bcd_in1=10010010 bcd_in2=01000110 cout=1 sum=00111000
* bcd_in1=10010010 bcd_in2=01000111 cout=1 sum=00111001
* bcd_in1=10010010 bcd_in2=01001000 cout=1 sum=01000000
* bcd_in1=10010010 bcd_in2=01001001 cout=1 sum=01000001
* bcd_in1=10010010 bcd_in2=01010000 cout=1 sum=01000010
* bcd_in1=10010010 bcd_in2=01010001 cout=1 sum=01000011
* bcd_in1=10010010 bcd_in2=01010010 cout=1 sum=01000100
* bcd_in1=10010010 bcd_in2=01010011 cout=1 sum=01000101
* bcd_in1=10010010 bcd_in2=01010100 cout=1 sum=01000110
* bcd_in1=10010010 bcd_in2=01010101 cout=1 sum=01000111
* bcd_in1=10010010 bcd_in2=01010110 cout=1 sum=01001000
* bcd_in1=10010010 bcd_in2=01010111 cout=1 sum=01001001
* bcd_in1=10010010 bcd_in2=01011000 cout=1 sum=01010000
* bcd_in1=10010010 bcd_in2=01011001 cout=1 sum=01010001
* bcd_in1=10010010 bcd_in2=01100000 cout=1 sum=01010010
* bcd_in1=10010010 bcd_in2=01100001 cout=1 sum=01010011
* bcd_in1=10010010 bcd_in2=01100010 cout=1 sum=01010100
* bcd_in1=10010010 bcd_in2=01100011 cout=1 sum=01010101
* bcd_in1=10010010 bcd_in2=01100100 cout=1 sum=01010110
* bcd_in1=10010010 bcd_in2=01100101 cout=1 sum=01010111
* bcd_in1=10010010 bcd_in2=01100110 cout=1 sum=01011000
* bcd_in1=10010010 bcd_in2=01100111 cout=1 sum=01011001
* bcd_in1=10010010 bcd_in2=01101000 cout=1 sum=01100000
* bcd_in1=10010010 bcd_in2=01101001 cout=1 sum=01100001
* bcd_in1=10010010 bcd_in2=01110000 cout=1 sum=01100010
* bcd_in1=10010010 bcd_in2=01110001 cout=1 sum=01100011
* bcd_in1=10010010 bcd_in2=01110010 cout=1 sum=01100100
* bcd_in1=10010010 bcd_in2=01110011 cout=1 sum=01100101
* bcd_in1=10010010 bcd_in2=01110100 cout=1 sum=01100110
* bcd_in1=10010010 bcd_in2=01110101 cout=1 sum=01100111
* bcd_in1=10010010 bcd_in2=01110110 cout=1 sum=01101000
* bcd_in1=10010010 bcd_in2=01110111 cout=1 sum=01101001
* bcd_in1=10010010 bcd_in2=01111000 cout=1 sum=01110000
* bcd_in1=10010010 bcd_in2=01111001 cout=1 sum=01110001
* bcd_in1=10010010 bcd_in2=10000000 cout=1 sum=01110010
* bcd_in1=10010010 bcd_in2=10000001 cout=1 sum=01110011
* bcd_in1=10010010 bcd_in2=10000010 cout=1 sum=01110100
* bcd_in1=10010010 bcd_in2=10000011 cout=1 sum=01110101
* bcd_in1=10010010 bcd_in2=10000100 cout=1 sum=01110110
* bcd_in1=10010010 bcd_in2=10000101 cout=1 sum=01110111
* bcd_in1=10010010 bcd_in2=10000110 cout=1 sum=01111000
* bcd_in1=10010010 bcd_in2=10000111 cout=1 sum=01111001
* bcd_in1=10010010 bcd_in2=10001000 cout=1 sum=10000000
* bcd_in1=10010010 bcd_in2=10001001 cout=1 sum=10000001
* bcd_in1=10010010 bcd_in2=10010000 cout=1 sum=10000010
* bcd_in1=10010010 bcd_in2=10010001 cout=1 sum=10000011
* bcd_in1=10010010 bcd_in2=10010010 cout=1 sum=10000100
* bcd_in1=10010010 bcd_in2=10010011 cout=1 sum=10000101
* bcd_in1=10010010 bcd_in2=10010100 cout=1 sum=10000110
* bcd_in1=10010010 bcd_in2=10010101 cout=1 sum=10000111
* bcd_in1=10010010 bcd_in2=10010110 cout=1 sum=10001000
* bcd_in1=10010010 bcd_in2=10010111 cout=1 sum=10001001
* bcd_in1=10010010 bcd_in2=10011000 cout=1 sum=10010000
* bcd_in1=10010010 bcd_in2=10011001 cout=1 sum=10010001
* bcd_in1=10010011 bcd_in2=00000000 cout=0 sum=10010011
* bcd_in1=10010011 bcd_in2=00000001 cout=0 sum=10010100
* bcd_in1=10010011 bcd_in2=00000010 cout=0 sum=10010101
* bcd_in1=10010011 bcd_in2=00000011 cout=0 sum=10010110
* bcd_in1=10010011 bcd_in2=00000100 cout=0 sum=10010111
* bcd_in1=10010011 bcd_in2=00000101 cout=0 sum=10011000
* bcd_in1=10010011 bcd_in2=00000110 cout=0 sum=10011001
* bcd_in1=10010011 bcd_in2=00000111 cout=1 sum=00000000
* bcd_in1=10010011 bcd_in2=00001000 cout=1 sum=00000001
* bcd_in1=10010011 bcd_in2=00001001 cout=1 sum=00000010
* bcd_in1=10010011 bcd_in2=00010000 cout=1 sum=00000011
* bcd_in1=10010011 bcd_in2=00010001 cout=1 sum=00000100
* bcd_in1=10010011 bcd_in2=00010010 cout=1 sum=00000101
* bcd_in1=10010011 bcd_in2=00010011 cout=1 sum=00000110
* bcd_in1=10010011 bcd_in2=00010100 cout=1 sum=00000111
* bcd_in1=10010011 bcd_in2=00010101 cout=1 sum=00001000
* bcd_in1=10010011 bcd_in2=00010110 cout=1 sum=00001001
* bcd_in1=10010011 bcd_in2=00010111 cout=1 sum=00010000
* bcd_in1=10010011 bcd_in2=00011000 cout=1 sum=00010001
* bcd_in1=10010011 bcd_in2=00011001 cout=1 sum=00010010
* bcd_in1=10010011 bcd_in2=00100000 cout=1 sum=00010011
* bcd_in1=10010011 bcd_in2=00100001 cout=1 sum=00010100
* bcd_in1=10010011 bcd_in2=00100010 cout=1 sum=00010101
* bcd_in1=10010011 bcd_in2=00100011 cout=1 sum=00010110
* bcd_in1=10010011 bcd_in2=00100100 cout=1 sum=00010111
* bcd_in1=10010011 bcd_in2=00100101 cout=1 sum=00011000
* bcd_in1=10010011 bcd_in2=00100110 cout=1 sum=00011001
* bcd_in1=10010011 bcd_in2=00100111 cout=1 sum=00100000
* bcd_in1=10010011 bcd_in2=00101000 cout=1 sum=00100001
* bcd_in1=10010011 bcd_in2=00101001 cout=1 sum=00100010
* bcd_in1=10010011 bcd_in2=00110000 cout=1 sum=00100011
* bcd_in1=10010011 bcd_in2=00110001 cout=1 sum=00100100
* bcd_in1=10010011 bcd_in2=00110010 cout=1 sum=00100101
* bcd_in1=10010011 bcd_in2=00110011 cout=1 sum=00100110
* bcd_in1=10010011 bcd_in2=00110100 cout=1 sum=00100111
* bcd_in1=10010011 bcd_in2=00110101 cout=1 sum=00101000
* bcd_in1=10010011 bcd_in2=00110110 cout=1 sum=00101001
* bcd_in1=10010011 bcd_in2=00110111 cout=1 sum=00110000
* bcd_in1=10010011 bcd_in2=00111000 cout=1 sum=00110001
* bcd_in1=10010011 bcd_in2=00111001 cout=1 sum=00110010
* bcd_in1=10010011 bcd_in2=01000000 cout=1 sum=00110011
* bcd_in1=10010011 bcd_in2=01000001 cout=1 sum=00110100
* bcd_in1=10010011 bcd_in2=01000010 cout=1 sum=00110101
* bcd_in1=10010011 bcd_in2=01000011 cout=1 sum=00110110
* bcd_in1=10010011 bcd_in2=01000100 cout=1 sum=00110111
* bcd_in1=10010011 bcd_in2=01000101 cout=1 sum=00111000
* bcd_in1=10010011 bcd_in2=01000110 cout=1 sum=00111001
* bcd_in1=10010011 bcd_in2=01000111 cout=1 sum=01000000
* bcd_in1=10010011 bcd_in2=01001000 cout=1 sum=01000001
* bcd_in1=10010011 bcd_in2=01001001 cout=1 sum=01000010
* bcd_in1=10010011 bcd_in2=01010000 cout=1 sum=01000011
* bcd_in1=10010011 bcd_in2=01010001 cout=1 sum=01000100
* bcd_in1=10010011 bcd_in2=01010010 cout=1 sum=01000101
* bcd_in1=10010011 bcd_in2=01010011 cout=1 sum=01000110
* bcd_in1=10010011 bcd_in2=01010100 cout=1 sum=01000111
* bcd_in1=10010011 bcd_in2=01010101 cout=1 sum=01001000
* bcd_in1=10010011 bcd_in2=01010110 cout=1 sum=01001001
* bcd_in1=10010011 bcd_in2=01010111 cout=1 sum=01010000
* bcd_in1=10010011 bcd_in2=01011000 cout=1 sum=01010001
* bcd_in1=10010011 bcd_in2=01011001 cout=1 sum=01010010
* bcd_in1=10010011 bcd_in2=01100000 cout=1 sum=01010011
* bcd_in1=10010011 bcd_in2=01100001 cout=1 sum=01010100
* bcd_in1=10010011 bcd_in2=01100010 cout=1 sum=01010101
* bcd_in1=10010011 bcd_in2=01100011 cout=1 sum=01010110
* bcd_in1=10010011 bcd_in2=01100100 cout=1 sum=01010111
* bcd_in1=10010011 bcd_in2=01100101 cout=1 sum=01011000
* bcd_in1=10010011 bcd_in2=01100110 cout=1 sum=01011001
* bcd_in1=10010011 bcd_in2=01100111 cout=1 sum=01100000
* bcd_in1=10010011 bcd_in2=01101000 cout=1 sum=01100001
* bcd_in1=10010011 bcd_in2=01101001 cout=1 sum=01100010
* bcd_in1=10010011 bcd_in2=01110000 cout=1 sum=01100011
* bcd_in1=10010011 bcd_in2=01110001 cout=1 sum=01100100
* bcd_in1=10010011 bcd_in2=01110010 cout=1 sum=01100101
* bcd_in1=10010011 bcd_in2=01110011 cout=1 sum=01100110
* bcd_in1=10010011 bcd_in2=01110100 cout=1 sum=01100111
* bcd_in1=10010011 bcd_in2=01110101 cout=1 sum=01101000
* bcd_in1=10010011 bcd_in2=01110110 cout=1 sum=01101001
* bcd_in1=10010011 bcd_in2=01110111 cout=1 sum=01110000
* bcd_in1=10010011 bcd_in2=01111000 cout=1 sum=01110001
* bcd_in1=10010011 bcd_in2=01111001 cout=1 sum=01110010
* bcd_in1=10010011 bcd_in2=10000000 cout=1 sum=01110011
* bcd_in1=10010011 bcd_in2=10000001 cout=1 sum=01110100
* bcd_in1=10010011 bcd_in2=10000010 cout=1 sum=01110101
* bcd_in1=10010011 bcd_in2=10000011 cout=1 sum=01110110
* bcd_in1=10010011 bcd_in2=10000100 cout=1 sum=01110111
* bcd_in1=10010011 bcd_in2=10000101 cout=1 sum=01111000
* bcd_in1=10010011 bcd_in2=10000110 cout=1 sum=01111001
* bcd_in1=10010011 bcd_in2=10000111 cout=1 sum=10000000
* bcd_in1=10010011 bcd_in2=10001000 cout=1 sum=10000001
* bcd_in1=10010011 bcd_in2=10001001 cout=1 sum=10000010
* bcd_in1=10010011 bcd_in2=10010000 cout=1 sum=10000011
* bcd_in1=10010011 bcd_in2=10010001 cout=1 sum=10000100
* bcd_in1=10010011 bcd_in2=10010010 cout=1 sum=10000101
* bcd_in1=10010011 bcd_in2=10010011 cout=1 sum=10000110
* bcd_in1=10010011 bcd_in2=10010100 cout=1 sum=10000111
* bcd_in1=10010011 bcd_in2=10010101 cout=1 sum=10001000
* bcd_in1=10010011 bcd_in2=10010110 cout=1 sum=10001001
* bcd_in1=10010011 bcd_in2=10010111 cout=1 sum=10010000
* bcd_in1=10010011 bcd_in2=10011000 cout=1 sum=10010001
* bcd_in1=10010011 bcd_in2=10011001 cout=1 sum=10010010
* bcd_in1=10010100 bcd_in2=00000000 cout=0 sum=10010100
* bcd_in1=10010100 bcd_in2=00000001 cout=0 sum=10010101
* bcd_in1=10010100 bcd_in2=00000010 cout=0 sum=10010110
* bcd_in1=10010100 bcd_in2=00000011 cout=0 sum=10010111
* bcd_in1=10010100 bcd_in2=00000100 cout=0 sum=10011000
* bcd_in1=10010100 bcd_in2=00000101 cout=0 sum=10011001
* bcd_in1=10010100 bcd_in2=00000110 cout=1 sum=00000000
* bcd_in1=10010100 bcd_in2=00000111 cout=1 sum=00000001
* bcd_in1=10010100 bcd_in2=00001000 cout=1 sum=00000010
* bcd_in1=10010100 bcd_in2=00001001 cout=1 sum=00000011
* bcd_in1=10010100 bcd_in2=00010000 cout=1 sum=00000100
* bcd_in1=10010100 bcd_in2=00010001 cout=1 sum=00000101
* bcd_in1=10010100 bcd_in2=00010010 cout=1 sum=00000110
* bcd_in1=10010100 bcd_in2=00010011 cout=1 sum=00000111
* bcd_in1=10010100 bcd_in2=00010100 cout=1 sum=00001000
* bcd_in1=10010100 bcd_in2=00010101 cout=1 sum=00001001
* bcd_in1=10010100 bcd_in2=00010110 cout=1 sum=00010000
* bcd_in1=10010100 bcd_in2=00010111 cout=1 sum=00010001
* bcd_in1=10010100 bcd_in2=00011000 cout=1 sum=00010010
* bcd_in1=10010100 bcd_in2=00011001 cout=1 sum=00010011
* bcd_in1=10010100 bcd_in2=00100000 cout=1 sum=00010100
* bcd_in1=10010100 bcd_in2=00100001 cout=1 sum=00010101
* bcd_in1=10010100 bcd_in2=00100010 cout=1 sum=00010110
* bcd_in1=10010100 bcd_in2=00100011 cout=1 sum=00010111
* bcd_in1=10010100 bcd_in2=00100100 cout=1 sum=00011000
* bcd_in1=10010100 bcd_in2=00100101 cout=1 sum=00011001
* bcd_in1=10010100 bcd_in2=00100110 cout=1 sum=00100000
* bcd_in1=10010100 bcd_in2=00100111 cout=1 sum=00100001
* bcd_in1=10010100 bcd_in2=00101000 cout=1 sum=00100010
* bcd_in1=10010100 bcd_in2=00101001 cout=1 sum=00100011
* bcd_in1=10010100 bcd_in2=00110000 cout=1 sum=00100100
* bcd_in1=10010100 bcd_in2=00110001 cout=1 sum=00100101
* bcd_in1=10010100 bcd_in2=00110010 cout=1 sum=00100110
* bcd_in1=10010100 bcd_in2=00110011 cout=1 sum=00100111
* bcd_in1=10010100 bcd_in2=00110100 cout=1 sum=00101000
* bcd_in1=10010100 bcd_in2=00110101 cout=1 sum=00101001
* bcd_in1=10010100 bcd_in2=00110110 cout=1 sum=00110000
* bcd_in1=10010100 bcd_in2=00110111 cout=1 sum=00110001
* bcd_in1=10010100 bcd_in2=00111000 cout=1 sum=00110010
* bcd_in1=10010100 bcd_in2=00111001 cout=1 sum=00110011
* bcd_in1=10010100 bcd_in2=01000000 cout=1 sum=00110100
* bcd_in1=10010100 bcd_in2=01000001 cout=1 sum=00110101
* bcd_in1=10010100 bcd_in2=01000010 cout=1 sum=00110110
* bcd_in1=10010100 bcd_in2=01000011 cout=1 sum=00110111
* bcd_in1=10010100 bcd_in2=01000100 cout=1 sum=00111000
* bcd_in1=10010100 bcd_in2=01000101 cout=1 sum=00111001
* bcd_in1=10010100 bcd_in2=01000110 cout=1 sum=01000000
* bcd_in1=10010100 bcd_in2=01000111 cout=1 sum=01000001
* bcd_in1=10010100 bcd_in2=01001000 cout=1 sum=01000010
* bcd_in1=10010100 bcd_in2=01001001 cout=1 sum=01000011
* bcd_in1=10010100 bcd_in2=01010000 cout=1 sum=01000100
* bcd_in1=10010100 bcd_in2=01010001 cout=1 sum=01000101
* bcd_in1=10010100 bcd_in2=01010010 cout=1 sum=01000110
* bcd_in1=10010100 bcd_in2=01010011 cout=1 sum=01000111
* bcd_in1=10010100 bcd_in2=01010100 cout=1 sum=01001000
* bcd_in1=10010100 bcd_in2=01010101 cout=1 sum=01001001
* bcd_in1=10010100 bcd_in2=01010110 cout=1 sum=01010000
* bcd_in1=10010100 bcd_in2=01010111 cout=1 sum=01010001
* bcd_in1=10010100 bcd_in2=01011000 cout=1 sum=01010010
* bcd_in1=10010100 bcd_in2=01011001 cout=1 sum=01010011
* bcd_in1=10010100 bcd_in2=01100000 cout=1 sum=01010100
* bcd_in1=10010100 bcd_in2=01100001 cout=1 sum=01010101
* bcd_in1=10010100 bcd_in2=01100010 cout=1 sum=01010110
* bcd_in1=10010100 bcd_in2=01100011 cout=1 sum=01010111
* bcd_in1=10010100 bcd_in2=01100100 cout=1 sum=01011000
* bcd_in1=10010100 bcd_in2=01100101 cout=1 sum=01011001
* bcd_in1=10010100 bcd_in2=01100110 cout=1 sum=01100000
* bcd_in1=10010100 bcd_in2=01100111 cout=1 sum=01100001
* bcd_in1=10010100 bcd_in2=01101000 cout=1 sum=01100010
* bcd_in1=10010100 bcd_in2=01101001 cout=1 sum=01100011
* bcd_in1=10010100 bcd_in2=01110000 cout=1 sum=01100100
* bcd_in1=10010100 bcd_in2=01110001 cout=1 sum=01100101
* bcd_in1=10010100 bcd_in2=01110010 cout=1 sum=01100110
* bcd_in1=10010100 bcd_in2=01110011 cout=1 sum=01100111
* bcd_in1=10010100 bcd_in2=01110100 cout=1 sum=01101000
* bcd_in1=10010100 bcd_in2=01110101 cout=1 sum=01101001
* bcd_in1=10010100 bcd_in2=01110110 cout=1 sum=01110000
* bcd_in1=10010100 bcd_in2=01110111 cout=1 sum=01110001
* bcd_in1=10010100 bcd_in2=01111000 cout=1 sum=01110010
* bcd_in1=10010100 bcd_in2=01111001 cout=1 sum=01110011
* bcd_in1=10010100 bcd_in2=10000000 cout=1 sum=01110100
* bcd_in1=10010100 bcd_in2=10000001 cout=1 sum=01110101
* bcd_in1=10010100 bcd_in2=10000010 cout=1 sum=01110110
* bcd_in1=10010100 bcd_in2=10000011 cout=1 sum=01110111
* bcd_in1=10010100 bcd_in2=10000100 cout=1 sum=01111000
* bcd_in1=10010100 bcd_in2=10000101 cout=1 sum=01111001
* bcd_in1=10010100 bcd_in2=10000110 cout=1 sum=10000000
* bcd_in1=10010100 bcd_in2=10000111 cout=1 sum=10000001
* bcd_in1=10010100 bcd_in2=10001000 cout=1 sum=10000010
* bcd_in1=10010100 bcd_in2=10001001 cout=1 sum=10000011
* bcd_in1=10010100 bcd_in2=10010000 cout=1 sum=10000100
* bcd_in1=10010100 bcd_in2=10010001 cout=1 sum=10000101
* bcd_in1=10010100 bcd_in2=10010010 cout=1 sum=10000110
* bcd_in1=10010100 bcd_in2=10010011 cout=1 sum=10000111
* bcd_in1=10010100 bcd_in2=10010100 cout=1 sum=10001000
* bcd_in1=10010100 bcd_in2=10010101 cout=1 sum=10001001
* bcd_in1=10010100 bcd_in2=10010110 cout=1 sum=10010000
* bcd_in1=10010100 bcd_in2=10010111 cout=1 sum=10010001
* bcd_in1=10010100 bcd_in2=10011000 cout=1 sum=10010010
* bcd_in1=10010100 bcd_in2=10011001 cout=1 sum=10010011
* bcd_in1=10010101 bcd_in2=00000000 cout=0 sum=10010101
* bcd_in1=10010101 bcd_in2=00000001 cout=0 sum=10010110
* bcd_in1=10010101 bcd_in2=00000010 cout=0 sum=10010111
* bcd_in1=10010101 bcd_in2=00000011 cout=0 sum=10011000
* bcd_in1=10010101 bcd_in2=00000100 cout=0 sum=10011001
* bcd_in1=10010101 bcd_in2=00000101 cout=1 sum=00000000
* bcd_in1=10010101 bcd_in2=00000110 cout=1 sum=00000001
* bcd_in1=10010101 bcd_in2=00000111 cout=1 sum=00000010
* bcd_in1=10010101 bcd_in2=00001000 cout=1 sum=00000011
* bcd_in1=10010101 bcd_in2=00001001 cout=1 sum=00000100
* bcd_in1=10010101 bcd_in2=00010000 cout=1 sum=00000101
* bcd_in1=10010101 bcd_in2=00010001 cout=1 sum=00000110
* bcd_in1=10010101 bcd_in2=00010010 cout=1 sum=00000111
* bcd_in1=10010101 bcd_in2=00010011 cout=1 sum=00001000
* bcd_in1=10010101 bcd_in2=00010100 cout=1 sum=00001001
* bcd_in1=10010101 bcd_in2=00010101 cout=1 sum=00010000
* bcd_in1=10010101 bcd_in2=00010110 cout=1 sum=00010001
* bcd_in1=10010101 bcd_in2=00010111 cout=1 sum=00010010
* bcd_in1=10010101 bcd_in2=00011000 cout=1 sum=00010011
* bcd_in1=10010101 bcd_in2=00011001 cout=1 sum=00010100
* bcd_in1=10010101 bcd_in2=00100000 cout=1 sum=00010101
* bcd_in1=10010101 bcd_in2=00100001 cout=1 sum=00010110
* bcd_in1=10010101 bcd_in2=00100010 cout=1 sum=00010111
* bcd_in1=10010101 bcd_in2=00100011 cout=1 sum=00011000
* bcd_in1=10010101 bcd_in2=00100100 cout=1 sum=00011001
* bcd_in1=10010101 bcd_in2=00100101 cout=1 sum=00100000
* bcd_in1=10010101 bcd_in2=00100110 cout=1 sum=00100001
* bcd_in1=10010101 bcd_in2=00100111 cout=1 sum=00100010
* bcd_in1=10010101 bcd_in2=00101000 cout=1 sum=00100011
* bcd_in1=10010101 bcd_in2=00101001 cout=1 sum=00100100
* bcd_in1=10010101 bcd_in2=00110000 cout=1 sum=00100101
* bcd_in1=10010101 bcd_in2=00110001 cout=1 sum=00100110
* bcd_in1=10010101 bcd_in2=00110010 cout=1 sum=00100111
* bcd_in1=10010101 bcd_in2=00110011 cout=1 sum=00101000
* bcd_in1=10010101 bcd_in2=00110100 cout=1 sum=00101001
* bcd_in1=10010101 bcd_in2=00110101 cout=1 sum=00110000
* bcd_in1=10010101 bcd_in2=00110110 cout=1 sum=00110001
* bcd_in1=10010101 bcd_in2=00110111 cout=1 sum=00110010
* bcd_in1=10010101 bcd_in2=00111000 cout=1 sum=00110011
* bcd_in1=10010101 bcd_in2=00111001 cout=1 sum=00110100
* bcd_in1=10010101 bcd_in2=01000000 cout=1 sum=00110101
* bcd_in1=10010101 bcd_in2=01000001 cout=1 sum=00110110
* bcd_in1=10010101 bcd_in2=01000010 cout=1 sum=00110111
* bcd_in1=10010101 bcd_in2=01000011 cout=1 sum=00111000
* bcd_in1=10010101 bcd_in2=01000100 cout=1 sum=00111001
* bcd_in1=10010101 bcd_in2=01000101 cout=1 sum=01000000
* bcd_in1=10010101 bcd_in2=01000110 cout=1 sum=01000001
* bcd_in1=10010101 bcd_in2=01000111 cout=1 sum=01000010
* bcd_in1=10010101 bcd_in2=01001000 cout=1 sum=01000011
* bcd_in1=10010101 bcd_in2=01001001 cout=1 sum=01000100
* bcd_in1=10010101 bcd_in2=01010000 cout=1 sum=01000101
* bcd_in1=10010101 bcd_in2=01010001 cout=1 sum=01000110
* bcd_in1=10010101 bcd_in2=01010010 cout=1 sum=01000111
* bcd_in1=10010101 bcd_in2=01010011 cout=1 sum=01001000
* bcd_in1=10010101 bcd_in2=01010100 cout=1 sum=01001001
* bcd_in1=10010101 bcd_in2=01010101 cout=1 sum=01010000
* bcd_in1=10010101 bcd_in2=01010110 cout=1 sum=01010001
* bcd_in1=10010101 bcd_in2=01010111 cout=1 sum=01010010
* bcd_in1=10010101 bcd_in2=01011000 cout=1 sum=01010011
* bcd_in1=10010101 bcd_in2=01011001 cout=1 sum=01010100
* bcd_in1=10010101 bcd_in2=01100000 cout=1 sum=01010101
* bcd_in1=10010101 bcd_in2=01100001 cout=1 sum=01010110
* bcd_in1=10010101 bcd_in2=01100010 cout=1 sum=01010111
* bcd_in1=10010101 bcd_in2=01100011 cout=1 sum=01011000
* bcd_in1=10010101 bcd_in2=01100100 cout=1 sum=01011001
* bcd_in1=10010101 bcd_in2=01100101 cout=1 sum=01100000
* bcd_in1=10010101 bcd_in2=01100110 cout=1 sum=01100001
* bcd_in1=10010101 bcd_in2=01100111 cout=1 sum=01100010
* bcd_in1=10010101 bcd_in2=01101000 cout=1 sum=01100011
* bcd_in1=10010101 bcd_in2=01101001 cout=1 sum=01100100
* bcd_in1=10010101 bcd_in2=01110000 cout=1 sum=01100101
* bcd_in1=10010101 bcd_in2=01110001 cout=1 sum=01100110
* bcd_in1=10010101 bcd_in2=01110010 cout=1 sum=01100111
* bcd_in1=10010101 bcd_in2=01110011 cout=1 sum=01101000
* bcd_in1=10010101 bcd_in2=01110100 cout=1 sum=01101001
* bcd_in1=10010101 bcd_in2=01110101 cout=1 sum=01110000
* bcd_in1=10010101 bcd_in2=01110110 cout=1 sum=01110001
* bcd_in1=10010101 bcd_in2=01110111 cout=1 sum=01110010
* bcd_in1=10010101 bcd_in2=01111000 cout=1 sum=01110011
* bcd_in1=10010101 bcd_in2=01111001 cout=1 sum=01110100
* bcd_in1=10010101 bcd_in2=10000000 cout=1 sum=01110101
* bcd_in1=10010101 bcd_in2=10000001 cout=1 sum=01110110
* bcd_in1=10010101 bcd_in2=10000010 cout=1 sum=01110111
* bcd_in1=10010101 bcd_in2=10000011 cout=1 sum=01111000
* bcd_in1=10010101 bcd_in2=10000100 cout=1 sum=01111001
* bcd_in1=10010101 bcd_in2=10000101 cout=1 sum=10000000
* bcd_in1=10010101 bcd_in2=10000110 cout=1 sum=10000001
* bcd_in1=10010101 bcd_in2=10000111 cout=1 sum=10000010
* bcd_in1=10010101 bcd_in2=10001000 cout=1 sum=10000011
* bcd_in1=10010101 bcd_in2=10001001 cout=1 sum=10000100
* bcd_in1=10010101 bcd_in2=10010000 cout=1 sum=10000101
* bcd_in1=10010101 bcd_in2=10010001 cout=1 sum=10000110
* bcd_in1=10010101 bcd_in2=10010010 cout=1 sum=10000111
* bcd_in1=10010101 bcd_in2=10010011 cout=1 sum=10001000
* bcd_in1=10010101 bcd_in2=10010100 cout=1 sum=10001001
* bcd_in1=10010101 bcd_in2=10010101 cout=1 sum=10010000
* bcd_in1=10010101 bcd_in2=10010110 cout=1 sum=10010001
* bcd_in1=10010101 bcd_in2=10010111 cout=1 sum=10010010
* bcd_in1=10010101 bcd_in2=10011000 cout=1 sum=10010011
* bcd_in1=10010101 bcd_in2=10011001 cout=1 sum=10010100
* bcd_in1=10010110 bcd_in2=00000000 cout=0 sum=10010110
* bcd_in1=10010110 bcd_in2=00000001 cout=0 sum=10010111
* bcd_in1=10010110 bcd_in2=00000010 cout=0 sum=10011000
* bcd_in1=10010110 bcd_in2=00000011 cout=0 sum=10011001
* bcd_in1=10010110 bcd_in2=00000100 cout=1 sum=00000000
* bcd_in1=10010110 bcd_in2=00000101 cout=1 sum=00000001
* bcd_in1=10010110 bcd_in2=00000110 cout=1 sum=00000010
* bcd_in1=10010110 bcd_in2=00000111 cout=1 sum=00000011
* bcd_in1=10010110 bcd_in2=00001000 cout=1 sum=00000100
* bcd_in1=10010110 bcd_in2=00001001 cout=1 sum=00000101
* bcd_in1=10010110 bcd_in2=00010000 cout=1 sum=00000110
* bcd_in1=10010110 bcd_in2=00010001 cout=1 sum=00000111
* bcd_in1=10010110 bcd_in2=00010010 cout=1 sum=00001000
* bcd_in1=10010110 bcd_in2=00010011 cout=1 sum=00001001
* bcd_in1=10010110 bcd_in2=00010100 cout=1 sum=00010000
* bcd_in1=10010110 bcd_in2=00010101 cout=1 sum=00010001
* bcd_in1=10010110 bcd_in2=00010110 cout=1 sum=00010010
* bcd_in1=10010110 bcd_in2=00010111 cout=1 sum=00010011
* bcd_in1=10010110 bcd_in2=00011000 cout=1 sum=00010100
* bcd_in1=10010110 bcd_in2=00011001 cout=1 sum=00010101
* bcd_in1=10010110 bcd_in2=00100000 cout=1 sum=00010110
* bcd_in1=10010110 bcd_in2=00100001 cout=1 sum=00010111
* bcd_in1=10010110 bcd_in2=00100010 cout=1 sum=00011000
* bcd_in1=10010110 bcd_in2=00100011 cout=1 sum=00011001
* bcd_in1=10010110 bcd_in2=00100100 cout=1 sum=00100000
* bcd_in1=10010110 bcd_in2=00100101 cout=1 sum=00100001
* bcd_in1=10010110 bcd_in2=00100110 cout=1 sum=00100010
* bcd_in1=10010110 bcd_in2=00100111 cout=1 sum=00100011
* bcd_in1=10010110 bcd_in2=00101000 cout=1 sum=00100100
* bcd_in1=10010110 bcd_in2=00101001 cout=1 sum=00100101
* bcd_in1=10010110 bcd_in2=00110000 cout=1 sum=00100110
* bcd_in1=10010110 bcd_in2=00110001 cout=1 sum=00100111
* bcd_in1=10010110 bcd_in2=00110010 cout=1 sum=00101000
* bcd_in1=10010110 bcd_in2=00110011 cout=1 sum=00101001
* bcd_in1=10010110 bcd_in2=00110100 cout=1 sum=00110000
* bcd_in1=10010110 bcd_in2=00110101 cout=1 sum=00110001
* bcd_in1=10010110 bcd_in2=00110110 cout=1 sum=00110010
* bcd_in1=10010110 bcd_in2=00110111 cout=1 sum=00110011
* bcd_in1=10010110 bcd_in2=00111000 cout=1 sum=00110100
* bcd_in1=10010110 bcd_in2=00111001 cout=1 sum=00110101
* bcd_in1=10010110 bcd_in2=01000000 cout=1 sum=00110110
* bcd_in1=10010110 bcd_in2=01000001 cout=1 sum=00110111
* bcd_in1=10010110 bcd_in2=01000010 cout=1 sum=00111000
* bcd_in1=10010110 bcd_in2=01000011 cout=1 sum=00111001
* bcd_in1=10010110 bcd_in2=01000100 cout=1 sum=01000000
* bcd_in1=10010110 bcd_in2=01000101 cout=1 sum=01000001
* bcd_in1=10010110 bcd_in2=01000110 cout=1 sum=01000010
* bcd_in1=10010110 bcd_in2=01000111 cout=1 sum=01000011
* bcd_in1=10010110 bcd_in2=01001000 cout=1 sum=01000100
* bcd_in1=10010110 bcd_in2=01001001 cout=1 sum=01000101
* bcd_in1=10010110 bcd_in2=01010000 cout=1 sum=01000110
* bcd_in1=10010110 bcd_in2=01010001 cout=1 sum=01000111
* bcd_in1=10010110 bcd_in2=01010010 cout=1 sum=01001000
* bcd_in1=10010110 bcd_in2=01010011 cout=1 sum=01001001
* bcd_in1=10010110 bcd_in2=01010100 cout=1 sum=01010000
* bcd_in1=10010110 bcd_in2=01010101 cout=1 sum=01010001
* bcd_in1=10010110 bcd_in2=01010110 cout=1 sum=01010010
* bcd_in1=10010110 bcd_in2=01010111 cout=1 sum=01010011
* bcd_in1=10010110 bcd_in2=01011000 cout=1 sum=01010100
* bcd_in1=10010110 bcd_in2=01011001 cout=1 sum=01010101
* bcd_in1=10010110 bcd_in2=01100000 cout=1 sum=01010110
* bcd_in1=10010110 bcd_in2=01100001 cout=1 sum=01010111
* bcd_in1=10010110 bcd_in2=01100010 cout=1 sum=01011000
* bcd_in1=10010110 bcd_in2=01100011 cout=1 sum=01011001
* bcd_in1=10010110 bcd_in2=01100100 cout=1 sum=01100000
* bcd_in1=10010110 bcd_in2=01100101 cout=1 sum=01100001
* bcd_in1=10010110 bcd_in2=01100110 cout=1 sum=01100010
* bcd_in1=10010110 bcd_in2=01100111 cout=1 sum=01100011
* bcd_in1=10010110 bcd_in2=01101000 cout=1 sum=01100100
* bcd_in1=10010110 bcd_in2=01101001 cout=1 sum=01100101
* bcd_in1=10010110 bcd_in2=01110000 cout=1 sum=01100110
* bcd_in1=10010110 bcd_in2=01110001 cout=1 sum=01100111
* bcd_in1=10010110 bcd_in2=01110010 cout=1 sum=01101000
* bcd_in1=10010110 bcd_in2=01110011 cout=1 sum=01101001
* bcd_in1=10010110 bcd_in2=01110100 cout=1 sum=01110000
* bcd_in1=10010110 bcd_in2=01110101 cout=1 sum=01110001
* bcd_in1=10010110 bcd_in2=01110110 cout=1 sum=01110010
* bcd_in1=10010110 bcd_in2=01110111 cout=1 sum=01110011
* bcd_in1=10010110 bcd_in2=01111000 cout=1 sum=01110100
* bcd_in1=10010110 bcd_in2=01111001 cout=1 sum=01110101
* bcd_in1=10010110 bcd_in2=10000000 cout=1 sum=01110110
* bcd_in1=10010110 bcd_in2=10000001 cout=1 sum=01110111
* bcd_in1=10010110 bcd_in2=10000010 cout=1 sum=01111000
* bcd_in1=10010110 bcd_in2=10000011 cout=1 sum=01111001
* bcd_in1=10010110 bcd_in2=10000100 cout=1 sum=10000000
* bcd_in1=10010110 bcd_in2=10000101 cout=1 sum=10000001
* bcd_in1=10010110 bcd_in2=10000110 cout=1 sum=10000010
* bcd_in1=10010110 bcd_in2=10000111 cout=1 sum=10000011
* bcd_in1=10010110 bcd_in2=10001000 cout=1 sum=10000100
* bcd_in1=10010110 bcd_in2=10001001 cout=1 sum=10000101
* bcd_in1=10010110 bcd_in2=10010000 cout=1 sum=10000110
* bcd_in1=10010110 bcd_in2=10010001 cout=1 sum=10000111
* bcd_in1=10010110 bcd_in2=10010010 cout=1 sum=10001000
* bcd_in1=10010110 bcd_in2=10010011 cout=1 sum=10001001
* bcd_in1=10010110 bcd_in2=10010100 cout=1 sum=10010000
* bcd_in1=10010110 bcd_in2=10010101 cout=1 sum=10010001
* bcd_in1=10010110 bcd_in2=10010110 cout=1 sum=10010010
* bcd_in1=10010110 bcd_in2=10010111 cout=1 sum=10010011
* bcd_in1=10010110 bcd_in2=10011000 cout=1 sum=10010100
* bcd_in1=10010110 bcd_in2=10011001 cout=1 sum=10010101
* bcd_in1=10010111 bcd_in2=00000000 cout=0 sum=10010111
* bcd_in1=10010111 bcd_in2=00000001 cout=0 sum=10011000
* bcd_in1=10010111 bcd_in2=00000010 cout=0 sum=10011001
* bcd_in1=10010111 bcd_in2=00000011 cout=1 sum=00000000
* bcd_in1=10010111 bcd_in2=00000100 cout=1 sum=00000001
* bcd_in1=10010111 bcd_in2=00000101 cout=1 sum=00000010
* bcd_in1=10010111 bcd_in2=00000110 cout=1 sum=00000011
* bcd_in1=10010111 bcd_in2=00000111 cout=1 sum=00000100
* bcd_in1=10010111 bcd_in2=00001000 cout=1 sum=00000101
* bcd_in1=10010111 bcd_in2=00001001 cout=1 sum=00000110
* bcd_in1=10010111 bcd_in2=00010000 cout=1 sum=00000111
* bcd_in1=10010111 bcd_in2=00010001 cout=1 sum=00001000
* bcd_in1=10010111 bcd_in2=00010010 cout=1 sum=00001001
* bcd_in1=10010111 bcd_in2=00010011 cout=1 sum=00010000
* bcd_in1=10010111 bcd_in2=00010100 cout=1 sum=00010001
* bcd_in1=10010111 bcd_in2=00010101 cout=1 sum=00010010
* bcd_in1=10010111 bcd_in2=00010110 cout=1 sum=00010011
* bcd_in1=10010111 bcd_in2=00010111 cout=1 sum=00010100
* bcd_in1=10010111 bcd_in2=00011000 cout=1 sum=00010101
* bcd_in1=10010111 bcd_in2=00011001 cout=1 sum=00010110
* bcd_in1=10010111 bcd_in2=00100000 cout=1 sum=00010111
* bcd_in1=10010111 bcd_in2=00100001 cout=1 sum=00011000
* bcd_in1=10010111 bcd_in2=00100010 cout=1 sum=00011001
* bcd_in1=10010111 bcd_in2=00100011 cout=1 sum=00100000
* bcd_in1=10010111 bcd_in2=00100100 cout=1 sum=00100001
* bcd_in1=10010111 bcd_in2=00100101 cout=1 sum=00100010
* bcd_in1=10010111 bcd_in2=00100110 cout=1 sum=00100011
* bcd_in1=10010111 bcd_in2=00100111 cout=1 sum=00100100
* bcd_in1=10010111 bcd_in2=00101000 cout=1 sum=00100101
* bcd_in1=10010111 bcd_in2=00101001 cout=1 sum=00100110
* bcd_in1=10010111 bcd_in2=00110000 cout=1 sum=00100111
* bcd_in1=10010111 bcd_in2=00110001 cout=1 sum=00101000
* bcd_in1=10010111 bcd_in2=00110010 cout=1 sum=00101001
* bcd_in1=10010111 bcd_in2=00110011 cout=1 sum=00110000
* bcd_in1=10010111 bcd_in2=00110100 cout=1 sum=00110001
* bcd_in1=10010111 bcd_in2=00110101 cout=1 sum=00110010
* bcd_in1=10010111 bcd_in2=00110110 cout=1 sum=00110011
* bcd_in1=10010111 bcd_in2=00110111 cout=1 sum=00110100
* bcd_in1=10010111 bcd_in2=00111000 cout=1 sum=00110101
* bcd_in1=10010111 bcd_in2=00111001 cout=1 sum=00110110
* bcd_in1=10010111 bcd_in2=01000000 cout=1 sum=00110111
* bcd_in1=10010111 bcd_in2=01000001 cout=1 sum=00111000
* bcd_in1=10010111 bcd_in2=01000010 cout=1 sum=00111001
* bcd_in1=10010111 bcd_in2=01000011 cout=1 sum=01000000
* bcd_in1=10010111 bcd_in2=01000100 cout=1 sum=01000001
* bcd_in1=10010111 bcd_in2=01000101 cout=1 sum=01000010
* bcd_in1=10010111 bcd_in2=01000110 cout=1 sum=01000011
* bcd_in1=10010111 bcd_in2=01000111 cout=1 sum=01000100
* bcd_in1=10010111 bcd_in2=01001000 cout=1 sum=01000101
* bcd_in1=10010111 bcd_in2=01001001 cout=1 sum=01000110
* bcd_in1=10010111 bcd_in2=01010000 cout=1 sum=01000111
* bcd_in1=10010111 bcd_in2=01010001 cout=1 sum=01001000
* bcd_in1=10010111 bcd_in2=01010010 cout=1 sum=01001001
* bcd_in1=10010111 bcd_in2=01010011 cout=1 sum=01010000
* bcd_in1=10010111 bcd_in2=01010100 cout=1 sum=01010001
* bcd_in1=10010111 bcd_in2=01010101 cout=1 sum=01010010
* bcd_in1=10010111 bcd_in2=01010110 cout=1 sum=01010011
* bcd_in1=10010111 bcd_in2=01010111 cout=1 sum=01010100
* bcd_in1=10010111 bcd_in2=01011000 cout=1 sum=01010101
* bcd_in1=10010111 bcd_in2=01011001 cout=1 sum=01010110
* bcd_in1=10010111 bcd_in2=01100000 cout=1 sum=01010111
* bcd_in1=10010111 bcd_in2=01100001 cout=1 sum=01011000
* bcd_in1=10010111 bcd_in2=01100010 cout=1 sum=01011001
* bcd_in1=10010111 bcd_in2=01100011 cout=1 sum=01100000
* bcd_in1=10010111 bcd_in2=01100100 cout=1 sum=01100001
* bcd_in1=10010111 bcd_in2=01100101 cout=1 sum=01100010
* bcd_in1=10010111 bcd_in2=01100110 cout=1 sum=01100011
* bcd_in1=10010111 bcd_in2=01100111 cout=1 sum=01100100
* bcd_in1=10010111 bcd_in2=01101000 cout=1 sum=01100101
* bcd_in1=10010111 bcd_in2=01101001 cout=1 sum=01100110
* bcd_in1=10010111 bcd_in2=01110000 cout=1 sum=01100111
* bcd_in1=10010111 bcd_in2=01110001 cout=1 sum=01101000
* bcd_in1=10010111 bcd_in2=01110010 cout=1 sum=01101001
* bcd_in1=10010111 bcd_in2=01110011 cout=1 sum=01110000
* bcd_in1=10010111 bcd_in2=01110100 cout=1 sum=01110001
* bcd_in1=10010111 bcd_in2=01110101 cout=1 sum=01110010
* bcd_in1=10010111 bcd_in2=01110110 cout=1 sum=01110011
* bcd_in1=10010111 bcd_in2=01110111 cout=1 sum=01110100
* bcd_in1=10010111 bcd_in2=01111000 cout=1 sum=01110101
* bcd_in1=10010111 bcd_in2=01111001 cout=1 sum=01110110
* bcd_in1=10010111 bcd_in2=10000000 cout=1 sum=01110111
* bcd_in1=10010111 bcd_in2=10000001 cout=1 sum=01111000
* bcd_in1=10010111 bcd_in2=10000010 cout=1 sum=01111001
* bcd_in1=10010111 bcd_in2=10000011 cout=1 sum=10000000
* bcd_in1=10010111 bcd_in2=10000100 cout=1 sum=10000001
* bcd_in1=10010111 bcd_in2=10000101 cout=1 sum=10000010
* bcd_in1=10010111 bcd_in2=10000110 cout=1 sum=10000011
* bcd_in1=10010111 bcd_in2=10000111 cout=1 sum=10000100
* bcd_in1=10010111 bcd_in2=10001000 cout=1 sum=10000101
* bcd_in1=10010111 bcd_in2=10001001 cout=1 sum=10000110
* bcd_in1=10010111 bcd_in2=10010000 cout=1 sum=10000111
* bcd_in1=10010111 bcd_in2=10010001 cout=1 sum=10001000
* bcd_in1=10010111 bcd_in2=10010010 cout=1 sum=10001001
* bcd_in1=10010111 bcd_in2=10010011 cout=1 sum=10010000
* bcd_in1=10010111 bcd_in2=10010100 cout=1 sum=10010001
* bcd_in1=10010111 bcd_in2=10010101 cout=1 sum=10010010
* bcd_in1=10010111 bcd_in2=10010110 cout=1 sum=10010011
* bcd_in1=10010111 bcd_in2=10010111 cout=1 sum=10010100
* bcd_in1=10010111 bcd_in2=10011000 cout=1 sum=10010101
* bcd_in1=10010111 bcd_in2=10011001 cout=1 sum=10010110
* bcd_in1=10011000 bcd_in2=00000000 cout=0 sum=10011000
* bcd_in1=10011000 bcd_in2=00000001 cout=0 sum=10011001
* bcd_in1=10011000 bcd_in2=00000010 cout=1 sum=00000000
* bcd_in1=10011000 bcd_in2=00000011 cout=1 sum=00000001
* bcd_in1=10011000 bcd_in2=00000100 cout=1 sum=00000010
* bcd_in1=10011000 bcd_in2=00000101 cout=1 sum=00000011
* bcd_in1=10011000 bcd_in2=00000110 cout=1 sum=00000100
* bcd_in1=10011000 bcd_in2=00000111 cout=1 sum=00000101
* bcd_in1=10011000 bcd_in2=00001000 cout=1 sum=00000110
* bcd_in1=10011000 bcd_in2=00001001 cout=1 sum=00000111
* bcd_in1=10011000 bcd_in2=00010000 cout=1 sum=00001000
* bcd_in1=10011000 bcd_in2=00010001 cout=1 sum=00001001
* bcd_in1=10011000 bcd_in2=00010010 cout=1 sum=00010000
* bcd_in1=10011000 bcd_in2=00010011 cout=1 sum=00010001
* bcd_in1=10011000 bcd_in2=00010100 cout=1 sum=00010010
* bcd_in1=10011000 bcd_in2=00010101 cout=1 sum=00010011
* bcd_in1=10011000 bcd_in2=00010110 cout=1 sum=00010100
* bcd_in1=10011000 bcd_in2=00010111 cout=1 sum=00010101
* bcd_in1=10011000 bcd_in2=00011000 cout=1 sum=00010110
* bcd_in1=10011000 bcd_in2=00011001 cout=1 sum=00010111
* bcd_in1=10011000 bcd_in2=00100000 cout=1 sum=00011000
* bcd_in1=10011000 bcd_in2=00100001 cout=1 sum=00011001
* bcd_in1=10011000 bcd_in2=00100010 cout=1 sum=00100000
* bcd_in1=10011000 bcd_in2=00100011 cout=1 sum=00100001
* bcd_in1=10011000 bcd_in2=00100100 cout=1 sum=00100010
* bcd_in1=10011000 bcd_in2=00100101 cout=1 sum=00100011
* bcd_in1=10011000 bcd_in2=00100110 cout=1 sum=00100100
* bcd_in1=10011000 bcd_in2=00100111 cout=1 sum=00100101
* bcd_in1=10011000 bcd_in2=00101000 cout=1 sum=00100110
* bcd_in1=10011000 bcd_in2=00101001 cout=1 sum=00100111
* bcd_in1=10011000 bcd_in2=00110000 cout=1 sum=00101000
* bcd_in1=10011000 bcd_in2=00110001 cout=1 sum=00101001
* bcd_in1=10011000 bcd_in2=00110010 cout=1 sum=00110000
* bcd_in1=10011000 bcd_in2=00110011 cout=1 sum=00110001
* bcd_in1=10011000 bcd_in2=00110100 cout=1 sum=00110010
* bcd_in1=10011000 bcd_in2=00110101 cout=1 sum=00110011
* bcd_in1=10011000 bcd_in2=00110110 cout=1 sum=00110100
* bcd_in1=10011000 bcd_in2=00110111 cout=1 sum=00110101
* bcd_in1=10011000 bcd_in2=00111000 cout=1 sum=00110110
* bcd_in1=10011000 bcd_in2=00111001 cout=1 sum=00110111
* bcd_in1=10011000 bcd_in2=01000000 cout=1 sum=00111000
* bcd_in1=10011000 bcd_in2=01000001 cout=1 sum=00111001
* bcd_in1=10011000 bcd_in2=01000010 cout=1 sum=01000000
* bcd_in1=10011000 bcd_in2=01000011 cout=1 sum=01000001
* bcd_in1=10011000 bcd_in2=01000100 cout=1 sum=01000010
* bcd_in1=10011000 bcd_in2=01000101 cout=1 sum=01000011
* bcd_in1=10011000 bcd_in2=01000110 cout=1 sum=01000100
* bcd_in1=10011000 bcd_in2=01000111 cout=1 sum=01000101
* bcd_in1=10011000 bcd_in2=01001000 cout=1 sum=01000110
* bcd_in1=10011000 bcd_in2=01001001 cout=1 sum=01000111
* bcd_in1=10011000 bcd_in2=01010000 cout=1 sum=01001000
* bcd_in1=10011000 bcd_in2=01010001 cout=1 sum=01001001
* bcd_in1=10011000 bcd_in2=01010010 cout=1 sum=01010000
* bcd_in1=10011000 bcd_in2=01010011 cout=1 sum=01010001
* bcd_in1=10011000 bcd_in2=01010100 cout=1 sum=01010010
* bcd_in1=10011000 bcd_in2=01010101 cout=1 sum=01010011
* bcd_in1=10011000 bcd_in2=01010110 cout=1 sum=01010100
* bcd_in1=10011000 bcd_in2=01010111 cout=1 sum=01010101
* bcd_in1=10011000 bcd_in2=01011000 cout=1 sum=01010110
* bcd_in1=10011000 bcd_in2=01011001 cout=1 sum=01010111
* bcd_in1=10011000 bcd_in2=01100000 cout=1 sum=01011000
* bcd_in1=10011000 bcd_in2=01100001 cout=1 sum=01011001
* bcd_in1=10011000 bcd_in2=01100010 cout=1 sum=01100000
* bcd_in1=10011000 bcd_in2=01100011 cout=1 sum=01100001
* bcd_in1=10011000 bcd_in2=01100100 cout=1 sum=01100010
* bcd_in1=10011000 bcd_in2=01100101 cout=1 sum=01100011
* bcd_in1=10011000 bcd_in2=01100110 cout=1 sum=01100100
* bcd_in1=10011000 bcd_in2=01100111 cout=1 sum=01100101
* bcd_in1=10011000 bcd_in2=01101000 cout=1 sum=01100110
* bcd_in1=10011000 bcd_in2=01101001 cout=1 sum=01100111
* bcd_in1=10011000 bcd_in2=01110000 cout=1 sum=01101000
* bcd_in1=10011000 bcd_in2=01110001 cout=1 sum=01101001
* bcd_in1=10011000 bcd_in2=01110010 cout=1 sum=01110000
* bcd_in1=10011000 bcd_in2=01110011 cout=1 sum=01110001
* bcd_in1=10011000 bcd_in2=01110100 cout=1 sum=01110010
* bcd_in1=10011000 bcd_in2=01110101 cout=1 sum=01110011
* bcd_in1=10011000 bcd_in2=01110110 cout=1 sum=01110100
* bcd_in1=10011000 bcd_in2=01110111 cout=1 sum=01110101
* bcd_in1=10011000 bcd_in2=01111000 cout=1 sum=01110110
* bcd_in1=10011000 bcd_in2=01111001 cout=1 sum=01110111
* bcd_in1=10011000 bcd_in2=10000000 cout=1 sum=01111000
* bcd_in1=10011000 bcd_in2=10000001 cout=1 sum=01111001
* bcd_in1=10011000 bcd_in2=10000010 cout=1 sum=10000000
* bcd_in1=10011000 bcd_in2=10000011 cout=1 sum=10000001
* bcd_in1=10011000 bcd_in2=10000100 cout=1 sum=10000010
* bcd_in1=10011000 bcd_in2=10000101 cout=1 sum=10000011
* bcd_in1=10011000 bcd_in2=10000110 cout=1 sum=10000100
* bcd_in1=10011000 bcd_in2=10000111 cout=1 sum=10000101
* bcd_in1=10011000 bcd_in2=10001000 cout=1 sum=10000110
* bcd_in1=10011000 bcd_in2=10001001 cout=1 sum=10000111
* bcd_in1=10011000 bcd_in2=10010000 cout=1 sum=10001000
* bcd_in1=10011000 bcd_in2=10010001 cout=1 sum=10001001
* bcd_in1=10011000 bcd_in2=10010010 cout=1 sum=10010000
* bcd_in1=10011000 bcd_in2=10010011 cout=1 sum=10010001
* bcd_in1=10011000 bcd_in2=10010100 cout=1 sum=10010010
* bcd_in1=10011000 bcd_in2=10010101 cout=1 sum=10010011
* bcd_in1=10011000 bcd_in2=10010110 cout=1 sum=10010100
* bcd_in1=10011000 bcd_in2=10010111 cout=1 sum=10010101
* bcd_in1=10011000 bcd_in2=10011000 cout=1 sum=10010110
* bcd_in1=10011000 bcd_in2=10011001 cout=1 sum=10010111
* bcd_in1=10011001 bcd_in2=00000000 cout=0 sum=10011001
* bcd_in1=10011001 bcd_in2=00000001 cout=1 sum=00000000
* bcd_in1=10011001 bcd_in2=00000010 cout=1 sum=00000001
* bcd_in1=10011001 bcd_in2=00000011 cout=1 sum=00000010
* bcd_in1=10011001 bcd_in2=00000100 cout=1 sum=00000011
* bcd_in1=10011001 bcd_in2=00000101 cout=1 sum=00000100
* bcd_in1=10011001 bcd_in2=00000110 cout=1 sum=00000101
* bcd_in1=10011001 bcd_in2=00000111 cout=1 sum=00000110
* bcd_in1=10011001 bcd_in2=00001000 cout=1 sum=00000111
* bcd_in1=10011001 bcd_in2=00001001 cout=1 sum=00001000
* bcd_in1=10011001 bcd_in2=00010000 cout=1 sum=00001001
* bcd_in1=10011001 bcd_in2=00010001 cout=1 sum=00010000
* bcd_in1=10011001 bcd_in2=00010010 cout=1 sum=00010001
* bcd_in1=10011001 bcd_in2=00010011 cout=1 sum=00010010
* bcd_in1=10011001 bcd_in2=00010100 cout=1 sum=00010011
* bcd_in1=10011001 bcd_in2=00010101 cout=1 sum=00010100
* bcd_in1=10011001 bcd_in2=00010110 cout=1 sum=00010101
* bcd_in1=10011001 bcd_in2=00010111 cout=1 sum=00010110
* bcd_in1=10011001 bcd_in2=00011000 cout=1 sum=00010111
* bcd_in1=10011001 bcd_in2=00011001 cout=1 sum=00011000
* bcd_in1=10011001 bcd_in2=00100000 cout=1 sum=00011001
* bcd_in1=10011001 bcd_in2=00100001 cout=1 sum=00100000
* bcd_in1=10011001 bcd_in2=00100010 cout=1 sum=00100001
* bcd_in1=10011001 bcd_in2=00100011 cout=1 sum=00100010
* bcd_in1=10011001 bcd_in2=00100100 cout=1 sum=00100011
* bcd_in1=10011001 bcd_in2=00100101 cout=1 sum=00100100
* bcd_in1=10011001 bcd_in2=00100110 cout=1 sum=00100101
* bcd_in1=10011001 bcd_in2=00100111 cout=1 sum=00100110
* bcd_in1=10011001 bcd_in2=00101000 cout=1 sum=00100111
* bcd_in1=10011001 bcd_in2=00101001 cout=1 sum=00101000
* bcd_in1=10011001 bcd_in2=00110000 cout=1 sum=00101001
* bcd_in1=10011001 bcd_in2=00110001 cout=1 sum=00110000
* bcd_in1=10011001 bcd_in2=00110010 cout=1 sum=00110001
* bcd_in1=10011001 bcd_in2=00110011 cout=1 sum=00110010
* bcd_in1=10011001 bcd_in2=00110100 cout=1 sum=00110011
* bcd_in1=10011001 bcd_in2=00110101 cout=1 sum=00110100
* bcd_in1=10011001 bcd_in2=00110110 cout=1 sum=00110101
* bcd_in1=10011001 bcd_in2=00110111 cout=1 sum=00110110
* bcd_in1=10011001 bcd_in2=00111000 cout=1 sum=00110111
* bcd_in1=10011001 bcd_in2=00111001 cout=1 sum=00111000
* bcd_in1=10011001 bcd_in2=01000000 cout=1 sum=00111001
* bcd_in1=10011001 bcd_in2=01000001 cout=1 sum=01000000
* bcd_in1=10011001 bcd_in2=01000010 cout=1 sum=01000001
* bcd_in1=10011001 bcd_in2=01000011 cout=1 sum=01000010
* bcd_in1=10011001 bcd_in2=01000100 cout=1 sum=01000011
* bcd_in1=10011001 bcd_in2=01000101 cout=1 sum=01000100
* bcd_in1=10011001 bcd_in2=01000110 cout=1 sum=01000101
* bcd_in1=10011001 bcd_in2=01000111 cout=1 sum=01000110
* bcd_in1=10011001 bcd_in2=01001000 cout=1 sum=01000111
* bcd_in1=10011001 bcd_in2=01001001 cout=1 sum=01001000
* bcd_in1=10011001 bcd_in2=01010000 cout=1 sum=01001001
* bcd_in1=10011001 bcd_in2=01010001 cout=1 sum=01010000
* bcd_in1=10011001 bcd_in2=01010010 cout=1 sum=01010001
* bcd_in1=10011001 bcd_in2=01010011 cout=1 sum=01010010
* bcd_in1=10011001 bcd_in2=01010100 cout=1 sum=01010011
* bcd_in1=10011001 bcd_in2=01010101 cout=1 sum=01010100
* bcd_in1=10011001 bcd_in2=01010110 cout=1 sum=01010101
* bcd_in1=10011001 bcd_in2=01010111 cout=1 sum=01010110
* bcd_in1=10011001 bcd_in2=01011000 cout=1 sum=01010111
* bcd_in1=10011001 bcd_in2=01011001 cout=1 sum=01011000
* bcd_in1=10011001 bcd_in2=01100000 cout=1 sum=01011001
* bcd_in1=10011001 bcd_in2=01100001 cout=1 sum=01100000
* bcd_in1=10011001 bcd_in2=01100010 cout=1 sum=01100001
* bcd_in1=10011001 bcd_in2=01100011 cout=1 sum=01100010
* bcd_in1=10011001 bcd_in2=01100100 cout=1 sum=01100011
* bcd_in1=10011001 bcd_in2=01100101 cout=1 sum=01100100
* bcd_in1=10011001 bcd_in2=01100110 cout=1 sum=01100101
* bcd_in1=10011001 bcd_in2=01100111 cout=1 sum=01100110
* bcd_in1=10011001 bcd_in2=01101000 cout=1 sum=01100111
* bcd_in1=10011001 bcd_in2=01101001 cout=1 sum=01101000
* bcd_in1=10011001 bcd_in2=01110000 cout=1 sum=01101001
* bcd_in1=10011001 bcd_in2=01110001 cout=1 sum=01110000
* bcd_in1=10011001 bcd_in2=01110010 cout=1 sum=01110001
* bcd_in1=10011001 bcd_in2=01110011 cout=1 sum=01110010
* bcd_in1=10011001 bcd_in2=01110100 cout=1 sum=01110011
* bcd_in1=10011001 bcd_in2=01110101 cout=1 sum=01110100
* bcd_in1=10011001 bcd_in2=01110110 cout=1 sum=01110101
* bcd_in1=10011001 bcd_in2=01110111 cout=1 sum=01110110
* bcd_in1=10011001 bcd_in2=01111000 cout=1 sum=01110111
* bcd_in1=10011001 bcd_in2=01111001 cout=1 sum=01111000
* bcd_in1=10011001 bcd_in2=10000000 cout=1 sum=01111001
* bcd_in1=10011001 bcd_in2=10000001 cout=1 sum=10000000
* bcd_in1=10011001 bcd_in2=10000010 cout=1 sum=10000001
* bcd_in1=10011001 bcd_in2=10000011 cout=1 sum=10000010
* bcd_in1=10011001 bcd_in2=10000100 cout=1 sum=10000011
* bcd_in1=10011001 bcd_in2=10000101 cout=1 sum=10000100
* bcd_in1=10011001 bcd_in2=10000110 cout=1 sum=10000101
* bcd_in1=10011001 bcd_in2=10000111 cout=1 sum=10000110
* bcd_in1=10011001 bcd_in2=10001000 cout=1 sum=10000111
* bcd_in1=10011001 bcd_in2=10001001 cout=1 sum=10001000
* bcd_in1=10011001 bcd_in2=10010000 cout=1 sum=10001001
* bcd_in1=10011001 bcd_in2=10010001 cout=1 sum=10010000
* bcd_in1=10011001 bcd_in2=10010010 cout=1 sum=10010001
* bcd_in1=10011001 bcd_in2=10010011 cout=1 sum=10010010
* bcd_in1=10011001 bcd_in2=10010100 cout=1 sum=10010011
* bcd_in1=10011001 bcd_in2=10010101 cout=1 sum=10010100
* bcd_in1=10011001 bcd_in2=10010110 cout=1 sum=10010101
* bcd_in1=10011001 bcd_in2=10010111 cout=1 sum=10010110
* bcd_in1=10011001 bcd_in2=10011000 cout=1 sum=10010111
* bcd_in1=10011001 bcd_in2=10011001 cout=1 sum=10011000
* n_bit_bcd_adder_tb.v:48: $finish called at 101000 (1s)
* 
*/
