module _4bit_comparator_tb;
reg [3:0]a,b;
wire greater,equal,lesser;
_4bit_comparator dut(a,b,greater,equal,lesser);
integer i,j;
initial begin
    for(i=0;i<=15;i=i+1) begin
        a=i;
        for(j=0;j<=15;j=j+1) begin
            b=j;
            #10 $display("a=%b b=%b a>b=%b a==b=%b a<b=%b",a,b,greater,equal,lesser);
        end
        b=0;
    end
    $finish;
end
endmodule

/*
* OUTPUT
a=0000 b=0000 a>b=0 a==b=1 a<b=0
a=0000 b=0001 a>b=0 a==b=0 a<b=1
a=0000 b=0010 a>b=0 a==b=0 a<b=1
a=0000 b=0011 a>b=0 a==b=0 a<b=1
a=0000 b=0100 a>b=0 a==b=0 a<b=1
a=0000 b=0101 a>b=0 a==b=0 a<b=1
a=0000 b=0110 a>b=0 a==b=0 a<b=1
a=0000 b=0111 a>b=0 a==b=0 a<b=1
a=0000 b=1000 a>b=0 a==b=0 a<b=1
a=0000 b=1001 a>b=0 a==b=0 a<b=1
a=0000 b=1010 a>b=0 a==b=0 a<b=1
a=0000 b=1011 a>b=0 a==b=0 a<b=1
a=0000 b=1100 a>b=0 a==b=0 a<b=1
a=0000 b=1101 a>b=0 a==b=0 a<b=1
a=0000 b=1110 a>b=0 a==b=0 a<b=1
a=0000 b=1111 a>b=0 a==b=0 a<b=1
a=0001 b=0000 a>b=1 a==b=0 a<b=0
a=0001 b=0001 a>b=0 a==b=1 a<b=0
a=0001 b=0010 a>b=0 a==b=0 a<b=1
a=0001 b=0011 a>b=0 a==b=0 a<b=1
a=0001 b=0100 a>b=0 a==b=0 a<b=1
a=0001 b=0101 a>b=0 a==b=0 a<b=1
a=0001 b=0110 a>b=0 a==b=0 a<b=1
a=0001 b=0111 a>b=0 a==b=0 a<b=1
a=0001 b=1000 a>b=0 a==b=0 a<b=1
a=0001 b=1001 a>b=0 a==b=0 a<b=1
a=0001 b=1010 a>b=0 a==b=0 a<b=1
a=0001 b=1011 a>b=0 a==b=0 a<b=1
a=0001 b=1100 a>b=0 a==b=0 a<b=1
a=0001 b=1101 a>b=0 a==b=0 a<b=1
a=0001 b=1110 a>b=0 a==b=0 a<b=1
a=0001 b=1111 a>b=0 a==b=0 a<b=1
a=0010 b=0000 a>b=1 a==b=0 a<b=0
a=0010 b=0001 a>b=1 a==b=0 a<b=0
a=0010 b=0010 a>b=0 a==b=1 a<b=0
a=0010 b=0011 a>b=0 a==b=0 a<b=1
a=0010 b=0100 a>b=0 a==b=0 a<b=1
a=0010 b=0101 a>b=0 a==b=0 a<b=1
a=0010 b=0110 a>b=0 a==b=0 a<b=1
a=0010 b=0111 a>b=0 a==b=0 a<b=1
a=0010 b=1000 a>b=0 a==b=0 a<b=1
a=0010 b=1001 a>b=0 a==b=0 a<b=1
a=0010 b=1010 a>b=0 a==b=0 a<b=1
a=0010 b=1011 a>b=0 a==b=0 a<b=1
a=0010 b=1100 a>b=0 a==b=0 a<b=1
a=0010 b=1101 a>b=0 a==b=0 a<b=1
a=0010 b=1110 a>b=0 a==b=0 a<b=1
a=0010 b=1111 a>b=0 a==b=0 a<b=1
a=0011 b=0000 a>b=1 a==b=0 a<b=0
a=0011 b=0001 a>b=1 a==b=0 a<b=0
a=0011 b=0010 a>b=1 a==b=0 a<b=0
a=0011 b=0011 a>b=0 a==b=1 a<b=0
a=0011 b=0100 a>b=0 a==b=0 a<b=1
a=0011 b=0101 a>b=0 a==b=0 a<b=1
a=0011 b=0110 a>b=0 a==b=0 a<b=1
a=0011 b=0111 a>b=0 a==b=0 a<b=1
a=0011 b=1000 a>b=0 a==b=0 a<b=1
a=0011 b=1001 a>b=0 a==b=0 a<b=1
a=0011 b=1010 a>b=0 a==b=0 a<b=1
a=0011 b=1011 a>b=0 a==b=0 a<b=1
a=0011 b=1100 a>b=0 a==b=0 a<b=1
a=0011 b=1101 a>b=0 a==b=0 a<b=1
a=0011 b=1110 a>b=0 a==b=0 a<b=1
a=0011 b=1111 a>b=0 a==b=0 a<b=1
a=0100 b=0000 a>b=1 a==b=0 a<b=0
a=0100 b=0001 a>b=1 a==b=0 a<b=0
a=0100 b=0010 a>b=1 a==b=0 a<b=0
a=0100 b=0011 a>b=1 a==b=0 a<b=0
a=0100 b=0100 a>b=0 a==b=1 a<b=0
a=0100 b=0101 a>b=0 a==b=0 a<b=1
a=0100 b=0110 a>b=0 a==b=0 a<b=1
a=0100 b=0111 a>b=0 a==b=0 a<b=1
a=0100 b=1000 a>b=0 a==b=0 a<b=1
a=0100 b=1001 a>b=0 a==b=0 a<b=1
a=0100 b=1010 a>b=0 a==b=0 a<b=1
a=0100 b=1011 a>b=0 a==b=0 a<b=1
a=0100 b=1100 a>b=0 a==b=0 a<b=1
a=0100 b=1101 a>b=0 a==b=0 a<b=1
a=0100 b=1110 a>b=0 a==b=0 a<b=1
a=0100 b=1111 a>b=0 a==b=0 a<b=1
a=0101 b=0000 a>b=1 a==b=0 a<b=0
a=0101 b=0001 a>b=1 a==b=0 a<b=0
a=0101 b=0010 a>b=1 a==b=0 a<b=0
a=0101 b=0011 a>b=1 a==b=0 a<b=0
a=0101 b=0100 a>b=1 a==b=0 a<b=0
a=0101 b=0101 a>b=0 a==b=1 a<b=0
a=0101 b=0110 a>b=0 a==b=0 a<b=1
a=0101 b=0111 a>b=0 a==b=0 a<b=1
a=0101 b=1000 a>b=0 a==b=0 a<b=1
a=0101 b=1001 a>b=0 a==b=0 a<b=1
a=0101 b=1010 a>b=0 a==b=0 a<b=1
a=0101 b=1011 a>b=0 a==b=0 a<b=1
a=0101 b=1100 a>b=0 a==b=0 a<b=1
a=0101 b=1101 a>b=0 a==b=0 a<b=1
a=0101 b=1110 a>b=0 a==b=0 a<b=1
a=0101 b=1111 a>b=0 a==b=0 a<b=1
a=0110 b=0000 a>b=1 a==b=0 a<b=0
a=0110 b=0001 a>b=1 a==b=0 a<b=0
a=0110 b=0010 a>b=1 a==b=0 a<b=0
a=0110 b=0011 a>b=1 a==b=0 a<b=0
a=0110 b=0100 a>b=1 a==b=0 a<b=0
a=0110 b=0101 a>b=1 a==b=0 a<b=0
a=0110 b=0110 a>b=0 a==b=1 a<b=0
a=0110 b=0111 a>b=0 a==b=0 a<b=1
a=0110 b=1000 a>b=0 a==b=0 a<b=1
a=0110 b=1001 a>b=0 a==b=0 a<b=1
a=0110 b=1010 a>b=0 a==b=0 a<b=1
a=0110 b=1011 a>b=0 a==b=0 a<b=1
a=0110 b=1100 a>b=0 a==b=0 a<b=1
a=0110 b=1101 a>b=0 a==b=0 a<b=1
a=0110 b=1110 a>b=0 a==b=0 a<b=1
a=0110 b=1111 a>b=0 a==b=0 a<b=1
a=0111 b=0000 a>b=1 a==b=0 a<b=0
a=0111 b=0001 a>b=1 a==b=0 a<b=0
a=0111 b=0010 a>b=1 a==b=0 a<b=0
a=0111 b=0011 a>b=1 a==b=0 a<b=0
a=0111 b=0100 a>b=1 a==b=0 a<b=0
a=0111 b=0101 a>b=1 a==b=0 a<b=0
a=0111 b=0110 a>b=1 a==b=0 a<b=0
a=0111 b=0111 a>b=0 a==b=1 a<b=0
a=0111 b=1000 a>b=0 a==b=0 a<b=1
a=0111 b=1001 a>b=0 a==b=0 a<b=1
a=0111 b=1010 a>b=0 a==b=0 a<b=1
a=0111 b=1011 a>b=0 a==b=0 a<b=1
a=0111 b=1100 a>b=0 a==b=0 a<b=1
a=0111 b=1101 a>b=0 a==b=0 a<b=1
a=0111 b=1110 a>b=0 a==b=0 a<b=1
a=0111 b=1111 a>b=0 a==b=0 a<b=1
a=1000 b=0000 a>b=1 a==b=0 a<b=0
a=1000 b=0001 a>b=1 a==b=0 a<b=0
a=1000 b=0010 a>b=1 a==b=0 a<b=0
a=1000 b=0011 a>b=1 a==b=0 a<b=0
a=1000 b=0100 a>b=1 a==b=0 a<b=0
a=1000 b=0101 a>b=1 a==b=0 a<b=0
a=1000 b=0110 a>b=1 a==b=0 a<b=0
a=1000 b=0111 a>b=1 a==b=0 a<b=0
a=1000 b=1000 a>b=0 a==b=1 a<b=0
a=1000 b=1001 a>b=0 a==b=0 a<b=1
a=1000 b=1010 a>b=0 a==b=0 a<b=1
a=1000 b=1011 a>b=0 a==b=0 a<b=1
a=1000 b=1100 a>b=0 a==b=0 a<b=1
a=1000 b=1101 a>b=0 a==b=0 a<b=1
a=1000 b=1110 a>b=0 a==b=0 a<b=1
a=1000 b=1111 a>b=0 a==b=0 a<b=1
a=1001 b=0000 a>b=1 a==b=0 a<b=0
a=1001 b=0001 a>b=1 a==b=0 a<b=0
a=1001 b=0010 a>b=1 a==b=0 a<b=0
a=1001 b=0011 a>b=1 a==b=0 a<b=0
a=1001 b=0100 a>b=1 a==b=0 a<b=0
a=1001 b=0101 a>b=1 a==b=0 a<b=0
a=1001 b=0110 a>b=1 a==b=0 a<b=0
a=1001 b=0111 a>b=1 a==b=0 a<b=0
a=1001 b=1000 a>b=1 a==b=0 a<b=0
a=1001 b=1001 a>b=0 a==b=1 a<b=0
a=1001 b=1010 a>b=0 a==b=0 a<b=1
a=1001 b=1011 a>b=0 a==b=0 a<b=1
a=1001 b=1100 a>b=0 a==b=0 a<b=1
a=1001 b=1101 a>b=0 a==b=0 a<b=1
a=1001 b=1110 a>b=0 a==b=0 a<b=1
a=1001 b=1111 a>b=0 a==b=0 a<b=1
a=1010 b=0000 a>b=1 a==b=0 a<b=0
a=1010 b=0001 a>b=1 a==b=0 a<b=0
a=1010 b=0010 a>b=1 a==b=0 a<b=0
a=1010 b=0011 a>b=1 a==b=0 a<b=0
a=1010 b=0100 a>b=1 a==b=0 a<b=0
a=1010 b=0101 a>b=1 a==b=0 a<b=0
a=1010 b=0110 a>b=1 a==b=0 a<b=0
a=1010 b=0111 a>b=1 a==b=0 a<b=0
a=1010 b=1000 a>b=1 a==b=0 a<b=0
a=1010 b=1001 a>b=1 a==b=0 a<b=0
a=1010 b=1010 a>b=0 a==b=1 a<b=0
a=1010 b=1011 a>b=0 a==b=0 a<b=1
a=1010 b=1100 a>b=0 a==b=0 a<b=1
a=1010 b=1101 a>b=0 a==b=0 a<b=1
a=1010 b=1110 a>b=0 a==b=0 a<b=1
a=1010 b=1111 a>b=0 a==b=0 a<b=1
a=1011 b=0000 a>b=1 a==b=0 a<b=0
a=1011 b=0001 a>b=1 a==b=0 a<b=0
a=1011 b=0010 a>b=1 a==b=0 a<b=0
a=1011 b=0011 a>b=1 a==b=0 a<b=0
a=1011 b=0100 a>b=1 a==b=0 a<b=0
a=1011 b=0101 a>b=1 a==b=0 a<b=0
a=1011 b=0110 a>b=1 a==b=0 a<b=0
a=1011 b=0111 a>b=1 a==b=0 a<b=0
a=1011 b=1000 a>b=1 a==b=0 a<b=0
a=1011 b=1001 a>b=1 a==b=0 a<b=0
a=1011 b=1010 a>b=1 a==b=0 a<b=0
a=1011 b=1011 a>b=0 a==b=1 a<b=0
a=1011 b=1100 a>b=0 a==b=0 a<b=1
a=1011 b=1101 a>b=0 a==b=0 a<b=1
a=1011 b=1110 a>b=0 a==b=0 a<b=1
a=1011 b=1111 a>b=0 a==b=0 a<b=1
a=1100 b=0000 a>b=1 a==b=0 a<b=0
a=1100 b=0001 a>b=1 a==b=0 a<b=0
a=1100 b=0010 a>b=1 a==b=0 a<b=0
a=1100 b=0011 a>b=1 a==b=0 a<b=0
a=1100 b=0100 a>b=1 a==b=0 a<b=0
a=1100 b=0101 a>b=1 a==b=0 a<b=0
a=1100 b=0110 a>b=1 a==b=0 a<b=0
a=1100 b=0111 a>b=1 a==b=0 a<b=0
a=1100 b=1000 a>b=1 a==b=0 a<b=0
a=1100 b=1001 a>b=1 a==b=0 a<b=0
a=1100 b=1010 a>b=1 a==b=0 a<b=0
a=1100 b=1011 a>b=1 a==b=0 a<b=0
a=1100 b=1100 a>b=0 a==b=1 a<b=0
a=1100 b=1101 a>b=0 a==b=0 a<b=1
a=1100 b=1110 a>b=0 a==b=0 a<b=1
a=1100 b=1111 a>b=0 a==b=0 a<b=1
a=1101 b=0000 a>b=1 a==b=0 a<b=0
a=1101 b=0001 a>b=1 a==b=0 a<b=0
a=1101 b=0010 a>b=1 a==b=0 a<b=0
a=1101 b=0011 a>b=1 a==b=0 a<b=0
a=1101 b=0100 a>b=1 a==b=0 a<b=0
a=1101 b=0101 a>b=1 a==b=0 a<b=0
a=1101 b=0110 a>b=1 a==b=0 a<b=0
a=1101 b=0111 a>b=1 a==b=0 a<b=0
a=1101 b=1000 a>b=1 a==b=0 a<b=0
a=1101 b=1001 a>b=1 a==b=0 a<b=0
a=1101 b=1010 a>b=1 a==b=0 a<b=0
a=1101 b=1011 a>b=1 a==b=0 a<b=0
a=1101 b=1100 a>b=1 a==b=0 a<b=0
a=1101 b=1101 a>b=0 a==b=1 a<b=0
a=1101 b=1110 a>b=0 a==b=0 a<b=1
a=1101 b=1111 a>b=0 a==b=0 a<b=1
a=1110 b=0000 a>b=1 a==b=0 a<b=0
a=1110 b=0001 a>b=1 a==b=0 a<b=0
a=1110 b=0010 a>b=1 a==b=0 a<b=0
a=1110 b=0011 a>b=1 a==b=0 a<b=0
a=1110 b=0100 a>b=1 a==b=0 a<b=0
a=1110 b=0101 a>b=1 a==b=0 a<b=0
a=1110 b=0110 a>b=1 a==b=0 a<b=0
a=1110 b=0111 a>b=1 a==b=0 a<b=0
a=1110 b=1000 a>b=1 a==b=0 a<b=0
a=1110 b=1001 a>b=1 a==b=0 a<b=0
a=1110 b=1010 a>b=1 a==b=0 a<b=0
a=1110 b=1011 a>b=1 a==b=0 a<b=0
a=1110 b=1100 a>b=1 a==b=0 a<b=0
a=1110 b=1101 a>b=1 a==b=0 a<b=0
a=1110 b=1110 a>b=0 a==b=1 a<b=0
a=1110 b=1111 a>b=0 a==b=0 a<b=1
a=1111 b=0000 a>b=1 a==b=0 a<b=0
a=1111 b=0001 a>b=1 a==b=0 a<b=0
a=1111 b=0010 a>b=1 a==b=0 a<b=0
a=1111 b=0011 a>b=1 a==b=0 a<b=0
a=1111 b=0100 a>b=1 a==b=0 a<b=0
a=1111 b=0101 a>b=1 a==b=0 a<b=0
a=1111 b=0110 a>b=1 a==b=0 a<b=0
a=1111 b=0111 a>b=1 a==b=0 a<b=0
a=1111 b=1000 a>b=1 a==b=0 a<b=0
a=1111 b=1001 a>b=1 a==b=0 a<b=0
a=1111 b=1010 a>b=1 a==b=0 a<b=0
a=1111 b=1011 a>b=1 a==b=0 a<b=0
a=1111 b=1100 a>b=1 a==b=0 a<b=0
a=1111 b=1101 a>b=1 a==b=0 a<b=0
a=1111 b=1110 a>b=1 a==b=0 a<b=0
a=1111 b=1111 a>b=0 a==b=1 a<b=0
_4bit_comparator_tb.v:15: $finish called at 2560 (1s)
* 
*/
