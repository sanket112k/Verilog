module n_bit_bcd_to_2421_tb;
parameter N=2;
parameter B=N*$clog2(10);
reg [N*4-1:0]bcd_in;
wire [N*4-1:0]_2421_out;
n_bit_bcd_to_2421 #(.N(N)) dut1(
    .bcd_in(bcd_in),
    ._2421_out(_2421_out)
);
integer i,j,k;
reg [B+N*4:0]shift_reg;
initial begin
    shift_reg=0;
    for(k=0;k<=(2**B)-1;k=k+1) begin
        shift_reg[B-1:0]=k;
        for(i=0;i<B;i=i+1) begin
            for(j=0;j<B;j=j+1) begin
                if(shift_reg[B+j*4 +: 4]>=5)
                    shift_reg[B+j*4 +: 4] = shift_reg[B+j*4 +: 4] + 3;
            end
            shift_reg=shift_reg<<1;
        end
        if(shift_reg[B+N*4]==1) $finish;
        bcd_in<=shift_reg[B+N*4-1:B];#10;
        shift_reg[B+N*4:B]<=0;
    end
    $finish;
end
initial begin
    $monitor("bcd_in=%b _2421_out=%b",bcd_in,_2421_out);
end
endmodule


/*
* OUTPUT
bcd_in=00000000 _2421_out=00000000
bcd_in=00000001 _2421_out=00000001
bcd_in=00000010 _2421_out=00000010
bcd_in=00000011 _2421_out=00000011
bcd_in=00000100 _2421_out=00000100
bcd_in=00000101 _2421_out=00001011
bcd_in=00000110 _2421_out=00001100
bcd_in=00000111 _2421_out=00001101
bcd_in=00001000 _2421_out=00001110
bcd_in=00001001 _2421_out=00001111
bcd_in=00010000 _2421_out=00010000
bcd_in=00010001 _2421_out=00010001
bcd_in=00010010 _2421_out=00010010
bcd_in=00010011 _2421_out=00010011
bcd_in=00010100 _2421_out=00010100
bcd_in=00010101 _2421_out=00011011
bcd_in=00010110 _2421_out=00011100
bcd_in=00010111 _2421_out=00011101
bcd_in=00011000 _2421_out=00011110
bcd_in=00011001 _2421_out=00011111
bcd_in=00100000 _2421_out=00100000
bcd_in=00100001 _2421_out=00100001
bcd_in=00100010 _2421_out=00100010
bcd_in=00100011 _2421_out=00100011
bcd_in=00100100 _2421_out=00100100
bcd_in=00100101 _2421_out=00101011
bcd_in=00100110 _2421_out=00101100
bcd_in=00100111 _2421_out=00101101
bcd_in=00101000 _2421_out=00101110
bcd_in=00101001 _2421_out=00101111
bcd_in=00110000 _2421_out=00110000
bcd_in=00110001 _2421_out=00110001
bcd_in=00110010 _2421_out=00110010
bcd_in=00110011 _2421_out=00110011
bcd_in=00110100 _2421_out=00110100
bcd_in=00110101 _2421_out=00111011
bcd_in=00110110 _2421_out=00111100
bcd_in=00110111 _2421_out=00111101
bcd_in=00111000 _2421_out=00111110
bcd_in=00111001 _2421_out=00111111
bcd_in=01000000 _2421_out=01000000
bcd_in=01000001 _2421_out=01000001
bcd_in=01000010 _2421_out=01000010
bcd_in=01000011 _2421_out=01000011
bcd_in=01000100 _2421_out=01000100
bcd_in=01000101 _2421_out=01001011
bcd_in=01000110 _2421_out=01001100
bcd_in=01000111 _2421_out=01001101
bcd_in=01001000 _2421_out=01001110
bcd_in=01001001 _2421_out=01001111
bcd_in=01010000 _2421_out=10110000
bcd_in=01010001 _2421_out=10110001
bcd_in=01010010 _2421_out=10110010
bcd_in=01010011 _2421_out=10110011
bcd_in=01010100 _2421_out=10110100
bcd_in=01010101 _2421_out=10111011
bcd_in=01010110 _2421_out=10111100
bcd_in=01010111 _2421_out=10111101
bcd_in=01011000 _2421_out=10111110
bcd_in=01011001 _2421_out=10111111
bcd_in=01100000 _2421_out=11000000
bcd_in=01100001 _2421_out=11000001
bcd_in=01100010 _2421_out=11000010
bcd_in=01100011 _2421_out=11000011
bcd_in=01100100 _2421_out=11000100
bcd_in=01100101 _2421_out=11001011
bcd_in=01100110 _2421_out=11001100
bcd_in=01100111 _2421_out=11001101
bcd_in=01101000 _2421_out=11001110
bcd_in=01101001 _2421_out=11001111
bcd_in=01110000 _2421_out=11010000
bcd_in=01110001 _2421_out=11010001
bcd_in=01110010 _2421_out=11010010
bcd_in=01110011 _2421_out=11010011
bcd_in=01110100 _2421_out=11010100
bcd_in=01110101 _2421_out=11011011
bcd_in=01110110 _2421_out=11011100
bcd_in=01110111 _2421_out=11011101
bcd_in=01111000 _2421_out=11011110
bcd_in=01111001 _2421_out=11011111
bcd_in=10000000 _2421_out=11100000
bcd_in=10000001 _2421_out=11100001
bcd_in=10000010 _2421_out=11100010
bcd_in=10000011 _2421_out=11100011
bcd_in=10000100 _2421_out=11100100
bcd_in=10000101 _2421_out=11101011
bcd_in=10000110 _2421_out=11101100
bcd_in=10000111 _2421_out=11101101
bcd_in=10001000 _2421_out=11101110
bcd_in=10001001 _2421_out=11101111
bcd_in=10010000 _2421_out=11110000
bcd_in=10010001 _2421_out=11110001
bcd_in=10010010 _2421_out=11110010
bcd_in=10010011 _2421_out=11110011
bcd_in=10010100 _2421_out=11110100
bcd_in=10010101 _2421_out=11111011
bcd_in=10010110 _2421_out=11111100
bcd_in=10010111 _2421_out=11111101
bcd_in=10011000 _2421_out=11111110
bcd_in=10011001 _2421_out=11111111
n_bit_bcd_to_2421_tb.v:23: $finish called at 1000 (1s)
*/
