module first(output a,b);
	assign a=1'b0;
	assign b=1'b1;
endmodule
