module module_name(
	input a,b,
	output y
);
	assign y=a&b;
endmodule
