module part_select(input [7:0]in, output [3:0]out1, output [3:0]out2);
	assign {out1,out2}=in;
endmodule
