module bit_select(input [7:0]in, output sign);
	assign sign=in[7];
endmodule
