module conditional_operators(input [3:0]in, output out);
assign out=in[0]? 1:0;
endmodule
