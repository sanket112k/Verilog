module half_subtractor(
    input a,b,
    output diff
);
assign diff=a-b;
endmodule
