module binary_to_bcd_tb;
parameter N=10;
parameter D=(N*30103)/100000 + 1;
reg [N-1:0]bin_in;
wire [D*4-1:0]bcd_out;
integer i;
binary_to_bcd #(
    .N(N), 
    .D(D)
) dut(
    .bin_in(bin_in),
    .bcd_out(bcd_out)
);
initial begin
    for(i=0;i<=(2**N)-1;i=i+1) begin
        bin_in=i;
        #10 $display("bin_in=%b bcd_out=%b",bin_in,bcd_out);

    end
    $finish;
end
endmodule

/*
* OUTPUT
bin_in=0000000000 bcd_out=0000000000000000
bin_in=0000000001 bcd_out=0000000000000001
bin_in=0000000010 bcd_out=0000000000000010
bin_in=0000000011 bcd_out=0000000000000011
bin_in=0000000100 bcd_out=0000000000000100
bin_in=0000000101 bcd_out=0000000000000101
bin_in=0000000110 bcd_out=0000000000000110
bin_in=0000000111 bcd_out=0000000000000111
bin_in=0000001000 bcd_out=0000000000001000
bin_in=0000001001 bcd_out=0000000000001001
bin_in=0000001010 bcd_out=0000000000010000
bin_in=0000001011 bcd_out=0000000000010001
bin_in=0000001100 bcd_out=0000000000010010
bin_in=0000001101 bcd_out=0000000000010011
bin_in=0000001110 bcd_out=0000000000010100
bin_in=0000001111 bcd_out=0000000000010101
bin_in=0000010000 bcd_out=0000000000010110
bin_in=0000010001 bcd_out=0000000000010111
bin_in=0000010010 bcd_out=0000000000011000
bin_in=0000010011 bcd_out=0000000000011001
bin_in=0000010100 bcd_out=0000000000100000
bin_in=0000010101 bcd_out=0000000000100001
bin_in=0000010110 bcd_out=0000000000100010
bin_in=0000010111 bcd_out=0000000000100011
bin_in=0000011000 bcd_out=0000000000100100
bin_in=0000011001 bcd_out=0000000000100101
bin_in=0000011010 bcd_out=0000000000100110
bin_in=0000011011 bcd_out=0000000000100111
bin_in=0000011100 bcd_out=0000000000101000
bin_in=0000011101 bcd_out=0000000000101001
bin_in=0000011110 bcd_out=0000000000110000
bin_in=0000011111 bcd_out=0000000000110001
bin_in=0000100000 bcd_out=0000000000110010
bin_in=0000100001 bcd_out=0000000000110011
bin_in=0000100010 bcd_out=0000000000110100
bin_in=0000100011 bcd_out=0000000000110101
bin_in=0000100100 bcd_out=0000000000110110
bin_in=0000100101 bcd_out=0000000000110111
bin_in=0000100110 bcd_out=0000000000111000
bin_in=0000100111 bcd_out=0000000000111001
bin_in=0000101000 bcd_out=0000000001000000
bin_in=0000101001 bcd_out=0000000001000001
bin_in=0000101010 bcd_out=0000000001000010
bin_in=0000101011 bcd_out=0000000001000011
bin_in=0000101100 bcd_out=0000000001000100
bin_in=0000101101 bcd_out=0000000001000101
bin_in=0000101110 bcd_out=0000000001000110
bin_in=0000101111 bcd_out=0000000001000111
bin_in=0000110000 bcd_out=0000000001001000
bin_in=0000110001 bcd_out=0000000001001001
bin_in=0000110010 bcd_out=0000000001010000
bin_in=0000110011 bcd_out=0000000001010001
bin_in=0000110100 bcd_out=0000000001010010
bin_in=0000110101 bcd_out=0000000001010011
bin_in=0000110110 bcd_out=0000000001010100
bin_in=0000110111 bcd_out=0000000001010101
bin_in=0000111000 bcd_out=0000000001010110
bin_in=0000111001 bcd_out=0000000001010111
bin_in=0000111010 bcd_out=0000000001011000
bin_in=0000111011 bcd_out=0000000001011001
bin_in=0000111100 bcd_out=0000000001100000
bin_in=0000111101 bcd_out=0000000001100001
bin_in=0000111110 bcd_out=0000000001100010
bin_in=0000111111 bcd_out=0000000001100011
bin_in=0001000000 bcd_out=0000000001100100
bin_in=0001000001 bcd_out=0000000001100101
bin_in=0001000010 bcd_out=0000000001100110
bin_in=0001000011 bcd_out=0000000001100111
bin_in=0001000100 bcd_out=0000000001101000
bin_in=0001000101 bcd_out=0000000001101001
bin_in=0001000110 bcd_out=0000000001110000
bin_in=0001000111 bcd_out=0000000001110001
bin_in=0001001000 bcd_out=0000000001110010
bin_in=0001001001 bcd_out=0000000001110011
bin_in=0001001010 bcd_out=0000000001110100
bin_in=0001001011 bcd_out=0000000001110101
bin_in=0001001100 bcd_out=0000000001110110
bin_in=0001001101 bcd_out=0000000001110111
bin_in=0001001110 bcd_out=0000000001111000
bin_in=0001001111 bcd_out=0000000001111001
bin_in=0001010000 bcd_out=0000000010000000
bin_in=0001010001 bcd_out=0000000010000001
bin_in=0001010010 bcd_out=0000000010000010
bin_in=0001010011 bcd_out=0000000010000011
bin_in=0001010100 bcd_out=0000000010000100
bin_in=0001010101 bcd_out=0000000010000101
bin_in=0001010110 bcd_out=0000000010000110
bin_in=0001010111 bcd_out=0000000010000111
bin_in=0001011000 bcd_out=0000000010001000
bin_in=0001011001 bcd_out=0000000010001001
bin_in=0001011010 bcd_out=0000000010010000
bin_in=0001011011 bcd_out=0000000010010001
bin_in=0001011100 bcd_out=0000000010010010
bin_in=0001011101 bcd_out=0000000010010011
bin_in=0001011110 bcd_out=0000000010010100
bin_in=0001011111 bcd_out=0000000010010101
bin_in=0001100000 bcd_out=0000000010010110
bin_in=0001100001 bcd_out=0000000010010111
bin_in=0001100010 bcd_out=0000000010011000
bin_in=0001100011 bcd_out=0000000010011001
bin_in=0001100100 bcd_out=0000000100000000
bin_in=0001100101 bcd_out=0000000100000001
bin_in=0001100110 bcd_out=0000000100000010
bin_in=0001100111 bcd_out=0000000100000011
bin_in=0001101000 bcd_out=0000000100000100
bin_in=0001101001 bcd_out=0000000100000101
bin_in=0001101010 bcd_out=0000000100000110
bin_in=0001101011 bcd_out=0000000100000111
bin_in=0001101100 bcd_out=0000000100001000
bin_in=0001101101 bcd_out=0000000100001001
bin_in=0001101110 bcd_out=0000000100010000
bin_in=0001101111 bcd_out=0000000100010001
bin_in=0001110000 bcd_out=0000000100010010
bin_in=0001110001 bcd_out=0000000100010011
bin_in=0001110010 bcd_out=0000000100010100
bin_in=0001110011 bcd_out=0000000100010101
bin_in=0001110100 bcd_out=0000000100010110
bin_in=0001110101 bcd_out=0000000100010111
bin_in=0001110110 bcd_out=0000000100011000
bin_in=0001110111 bcd_out=0000000100011001
bin_in=0001111000 bcd_out=0000000100100000
bin_in=0001111001 bcd_out=0000000100100001
bin_in=0001111010 bcd_out=0000000100100010
bin_in=0001111011 bcd_out=0000000100100011
bin_in=0001111100 bcd_out=0000000100100100
bin_in=0001111101 bcd_out=0000000100100101
bin_in=0001111110 bcd_out=0000000100100110
bin_in=0001111111 bcd_out=0000000100100111
bin_in=0010000000 bcd_out=0000000100101000
bin_in=0010000001 bcd_out=0000000100101001
bin_in=0010000010 bcd_out=0000000100110000
bin_in=0010000011 bcd_out=0000000100110001
bin_in=0010000100 bcd_out=0000000100110010
bin_in=0010000101 bcd_out=0000000100110011
bin_in=0010000110 bcd_out=0000000100110100
bin_in=0010000111 bcd_out=0000000100110101
bin_in=0010001000 bcd_out=0000000100110110
bin_in=0010001001 bcd_out=0000000100110111
bin_in=0010001010 bcd_out=0000000100111000
bin_in=0010001011 bcd_out=0000000100111001
bin_in=0010001100 bcd_out=0000000101000000
bin_in=0010001101 bcd_out=0000000101000001
bin_in=0010001110 bcd_out=0000000101000010
bin_in=0010001111 bcd_out=0000000101000011
bin_in=0010010000 bcd_out=0000000101000100
bin_in=0010010001 bcd_out=0000000101000101
bin_in=0010010010 bcd_out=0000000101000110
bin_in=0010010011 bcd_out=0000000101000111
bin_in=0010010100 bcd_out=0000000101001000
bin_in=0010010101 bcd_out=0000000101001001
bin_in=0010010110 bcd_out=0000000101010000
bin_in=0010010111 bcd_out=0000000101010001
bin_in=0010011000 bcd_out=0000000101010010
bin_in=0010011001 bcd_out=0000000101010011
bin_in=0010011010 bcd_out=0000000101010100
bin_in=0010011011 bcd_out=0000000101010101
bin_in=0010011100 bcd_out=0000000101010110
bin_in=0010011101 bcd_out=0000000101010111
bin_in=0010011110 bcd_out=0000000101011000
bin_in=0010011111 bcd_out=0000000101011001
bin_in=0010100000 bcd_out=0000000101100000
bin_in=0010100001 bcd_out=0000000101100001
bin_in=0010100010 bcd_out=0000000101100010
bin_in=0010100011 bcd_out=0000000101100011
bin_in=0010100100 bcd_out=0000000101100100
bin_in=0010100101 bcd_out=0000000101100101
bin_in=0010100110 bcd_out=0000000101100110
bin_in=0010100111 bcd_out=0000000101100111
bin_in=0010101000 bcd_out=0000000101101000
bin_in=0010101001 bcd_out=0000000101101001
bin_in=0010101010 bcd_out=0000000101110000
bin_in=0010101011 bcd_out=0000000101110001
bin_in=0010101100 bcd_out=0000000101110010
bin_in=0010101101 bcd_out=0000000101110011
bin_in=0010101110 bcd_out=0000000101110100
bin_in=0010101111 bcd_out=0000000101110101
bin_in=0010110000 bcd_out=0000000101110110
bin_in=0010110001 bcd_out=0000000101110111
bin_in=0010110010 bcd_out=0000000101111000
bin_in=0010110011 bcd_out=0000000101111001
bin_in=0010110100 bcd_out=0000000110000000
bin_in=0010110101 bcd_out=0000000110000001
bin_in=0010110110 bcd_out=0000000110000010
bin_in=0010110111 bcd_out=0000000110000011
bin_in=0010111000 bcd_out=0000000110000100
bin_in=0010111001 bcd_out=0000000110000101
bin_in=0010111010 bcd_out=0000000110000110
bin_in=0010111011 bcd_out=0000000110000111
bin_in=0010111100 bcd_out=0000000110001000
bin_in=0010111101 bcd_out=0000000110001001
bin_in=0010111110 bcd_out=0000000110010000
bin_in=0010111111 bcd_out=0000000110010001
bin_in=0011000000 bcd_out=0000000110010010
bin_in=0011000001 bcd_out=0000000110010011
bin_in=0011000010 bcd_out=0000000110010100
bin_in=0011000011 bcd_out=0000000110010101
bin_in=0011000100 bcd_out=0000000110010110
bin_in=0011000101 bcd_out=0000000110010111
bin_in=0011000110 bcd_out=0000000110011000
bin_in=0011000111 bcd_out=0000000110011001
bin_in=0011001000 bcd_out=0000001000000000
bin_in=0011001001 bcd_out=0000001000000001
bin_in=0011001010 bcd_out=0000001000000010
bin_in=0011001011 bcd_out=0000001000000011
bin_in=0011001100 bcd_out=0000001000000100
bin_in=0011001101 bcd_out=0000001000000101
bin_in=0011001110 bcd_out=0000001000000110
bin_in=0011001111 bcd_out=0000001000000111
bin_in=0011010000 bcd_out=0000001000001000
bin_in=0011010001 bcd_out=0000001000001001
bin_in=0011010010 bcd_out=0000001000010000
bin_in=0011010011 bcd_out=0000001000010001
bin_in=0011010100 bcd_out=0000001000010010
bin_in=0011010101 bcd_out=0000001000010011
bin_in=0011010110 bcd_out=0000001000010100
bin_in=0011010111 bcd_out=0000001000010101
bin_in=0011011000 bcd_out=0000001000010110
bin_in=0011011001 bcd_out=0000001000010111
bin_in=0011011010 bcd_out=0000001000011000
bin_in=0011011011 bcd_out=0000001000011001
bin_in=0011011100 bcd_out=0000001000100000
bin_in=0011011101 bcd_out=0000001000100001
bin_in=0011011110 bcd_out=0000001000100010
bin_in=0011011111 bcd_out=0000001000100011
bin_in=0011100000 bcd_out=0000001000100100
bin_in=0011100001 bcd_out=0000001000100101
bin_in=0011100010 bcd_out=0000001000100110
bin_in=0011100011 bcd_out=0000001000100111
bin_in=0011100100 bcd_out=0000001000101000
bin_in=0011100101 bcd_out=0000001000101001
bin_in=0011100110 bcd_out=0000001000110000
bin_in=0011100111 bcd_out=0000001000110001
bin_in=0011101000 bcd_out=0000001000110010
bin_in=0011101001 bcd_out=0000001000110011
bin_in=0011101010 bcd_out=0000001000110100
bin_in=0011101011 bcd_out=0000001000110101
bin_in=0011101100 bcd_out=0000001000110110
bin_in=0011101101 bcd_out=0000001000110111
bin_in=0011101110 bcd_out=0000001000111000
bin_in=0011101111 bcd_out=0000001000111001
bin_in=0011110000 bcd_out=0000001001000000
bin_in=0011110001 bcd_out=0000001001000001
bin_in=0011110010 bcd_out=0000001001000010
bin_in=0011110011 bcd_out=0000001001000011
bin_in=0011110100 bcd_out=0000001001000100
bin_in=0011110101 bcd_out=0000001001000101
bin_in=0011110110 bcd_out=0000001001000110
bin_in=0011110111 bcd_out=0000001001000111
bin_in=0011111000 bcd_out=0000001001001000
bin_in=0011111001 bcd_out=0000001001001001
bin_in=0011111010 bcd_out=0000001001010000
bin_in=0011111011 bcd_out=0000001001010001
bin_in=0011111100 bcd_out=0000001001010010
bin_in=0011111101 bcd_out=0000001001010011
bin_in=0011111110 bcd_out=0000001001010100
bin_in=0011111111 bcd_out=0000001001010101
bin_in=0100000000 bcd_out=0000001001010110
bin_in=0100000001 bcd_out=0000001001010111
bin_in=0100000010 bcd_out=0000001001011000
bin_in=0100000011 bcd_out=0000001001011001
bin_in=0100000100 bcd_out=0000001001100000
bin_in=0100000101 bcd_out=0000001001100001
bin_in=0100000110 bcd_out=0000001001100010
bin_in=0100000111 bcd_out=0000001001100011
bin_in=0100001000 bcd_out=0000001001100100
bin_in=0100001001 bcd_out=0000001001100101
bin_in=0100001010 bcd_out=0000001001100110
bin_in=0100001011 bcd_out=0000001001100111
bin_in=0100001100 bcd_out=0000001001101000
bin_in=0100001101 bcd_out=0000001001101001
bin_in=0100001110 bcd_out=0000001001110000
bin_in=0100001111 bcd_out=0000001001110001
bin_in=0100010000 bcd_out=0000001001110010
bin_in=0100010001 bcd_out=0000001001110011
bin_in=0100010010 bcd_out=0000001001110100
bin_in=0100010011 bcd_out=0000001001110101
bin_in=0100010100 bcd_out=0000001001110110
bin_in=0100010101 bcd_out=0000001001110111
bin_in=0100010110 bcd_out=0000001001111000
bin_in=0100010111 bcd_out=0000001001111001
bin_in=0100011000 bcd_out=0000001010000000
bin_in=0100011001 bcd_out=0000001010000001
bin_in=0100011010 bcd_out=0000001010000010
bin_in=0100011011 bcd_out=0000001010000011
bin_in=0100011100 bcd_out=0000001010000100
bin_in=0100011101 bcd_out=0000001010000101
bin_in=0100011110 bcd_out=0000001010000110
bin_in=0100011111 bcd_out=0000001010000111
bin_in=0100100000 bcd_out=0000001010001000
bin_in=0100100001 bcd_out=0000001010001001
bin_in=0100100010 bcd_out=0000001010010000
bin_in=0100100011 bcd_out=0000001010010001
bin_in=0100100100 bcd_out=0000001010010010
bin_in=0100100101 bcd_out=0000001010010011
bin_in=0100100110 bcd_out=0000001010010100
bin_in=0100100111 bcd_out=0000001010010101
bin_in=0100101000 bcd_out=0000001010010110
bin_in=0100101001 bcd_out=0000001010010111
bin_in=0100101010 bcd_out=0000001010011000
bin_in=0100101011 bcd_out=0000001010011001
bin_in=0100101100 bcd_out=0000001100000000
bin_in=0100101101 bcd_out=0000001100000001
bin_in=0100101110 bcd_out=0000001100000010
bin_in=0100101111 bcd_out=0000001100000011
bin_in=0100110000 bcd_out=0000001100000100
bin_in=0100110001 bcd_out=0000001100000101
bin_in=0100110010 bcd_out=0000001100000110
bin_in=0100110011 bcd_out=0000001100000111
bin_in=0100110100 bcd_out=0000001100001000
bin_in=0100110101 bcd_out=0000001100001001
bin_in=0100110110 bcd_out=0000001100010000
bin_in=0100110111 bcd_out=0000001100010001
bin_in=0100111000 bcd_out=0000001100010010
bin_in=0100111001 bcd_out=0000001100010011
bin_in=0100111010 bcd_out=0000001100010100
bin_in=0100111011 bcd_out=0000001100010101
bin_in=0100111100 bcd_out=0000001100010110
bin_in=0100111101 bcd_out=0000001100010111
bin_in=0100111110 bcd_out=0000001100011000
bin_in=0100111111 bcd_out=0000001100011001
bin_in=0101000000 bcd_out=0000001100100000
bin_in=0101000001 bcd_out=0000001100100001
bin_in=0101000010 bcd_out=0000001100100010
bin_in=0101000011 bcd_out=0000001100100011
bin_in=0101000100 bcd_out=0000001100100100
bin_in=0101000101 bcd_out=0000001100100101
bin_in=0101000110 bcd_out=0000001100100110
bin_in=0101000111 bcd_out=0000001100100111
bin_in=0101001000 bcd_out=0000001100101000
bin_in=0101001001 bcd_out=0000001100101001
bin_in=0101001010 bcd_out=0000001100110000
bin_in=0101001011 bcd_out=0000001100110001
bin_in=0101001100 bcd_out=0000001100110010
bin_in=0101001101 bcd_out=0000001100110011
bin_in=0101001110 bcd_out=0000001100110100
bin_in=0101001111 bcd_out=0000001100110101
bin_in=0101010000 bcd_out=0000001100110110
bin_in=0101010001 bcd_out=0000001100110111
bin_in=0101010010 bcd_out=0000001100111000
bin_in=0101010011 bcd_out=0000001100111001
bin_in=0101010100 bcd_out=0000001101000000
bin_in=0101010101 bcd_out=0000001101000001
bin_in=0101010110 bcd_out=0000001101000010
bin_in=0101010111 bcd_out=0000001101000011
bin_in=0101011000 bcd_out=0000001101000100
bin_in=0101011001 bcd_out=0000001101000101
bin_in=0101011010 bcd_out=0000001101000110
bin_in=0101011011 bcd_out=0000001101000111
bin_in=0101011100 bcd_out=0000001101001000
bin_in=0101011101 bcd_out=0000001101001001
bin_in=0101011110 bcd_out=0000001101010000
bin_in=0101011111 bcd_out=0000001101010001
bin_in=0101100000 bcd_out=0000001101010010
bin_in=0101100001 bcd_out=0000001101010011
bin_in=0101100010 bcd_out=0000001101010100
bin_in=0101100011 bcd_out=0000001101010101
bin_in=0101100100 bcd_out=0000001101010110
bin_in=0101100101 bcd_out=0000001101010111
bin_in=0101100110 bcd_out=0000001101011000
bin_in=0101100111 bcd_out=0000001101011001
bin_in=0101101000 bcd_out=0000001101100000
bin_in=0101101001 bcd_out=0000001101100001
bin_in=0101101010 bcd_out=0000001101100010
bin_in=0101101011 bcd_out=0000001101100011
bin_in=0101101100 bcd_out=0000001101100100
bin_in=0101101101 bcd_out=0000001101100101
bin_in=0101101110 bcd_out=0000001101100110
bin_in=0101101111 bcd_out=0000001101100111
bin_in=0101110000 bcd_out=0000001101101000
bin_in=0101110001 bcd_out=0000001101101001
bin_in=0101110010 bcd_out=0000001101110000
bin_in=0101110011 bcd_out=0000001101110001
bin_in=0101110100 bcd_out=0000001101110010
bin_in=0101110101 bcd_out=0000001101110011
bin_in=0101110110 bcd_out=0000001101110100
bin_in=0101110111 bcd_out=0000001101110101
bin_in=0101111000 bcd_out=0000001101110110
bin_in=0101111001 bcd_out=0000001101110111
bin_in=0101111010 bcd_out=0000001101111000
bin_in=0101111011 bcd_out=0000001101111001
bin_in=0101111100 bcd_out=0000001110000000
bin_in=0101111101 bcd_out=0000001110000001
bin_in=0101111110 bcd_out=0000001110000010
bin_in=0101111111 bcd_out=0000001110000011
bin_in=0110000000 bcd_out=0000001110000100
bin_in=0110000001 bcd_out=0000001110000101
bin_in=0110000010 bcd_out=0000001110000110
bin_in=0110000011 bcd_out=0000001110000111
bin_in=0110000100 bcd_out=0000001110001000
bin_in=0110000101 bcd_out=0000001110001001
bin_in=0110000110 bcd_out=0000001110010000
bin_in=0110000111 bcd_out=0000001110010001
bin_in=0110001000 bcd_out=0000001110010010
bin_in=0110001001 bcd_out=0000001110010011
bin_in=0110001010 bcd_out=0000001110010100
bin_in=0110001011 bcd_out=0000001110010101
bin_in=0110001100 bcd_out=0000001110010110
bin_in=0110001101 bcd_out=0000001110010111
bin_in=0110001110 bcd_out=0000001110011000
bin_in=0110001111 bcd_out=0000001110011001
bin_in=0110010000 bcd_out=0000010000000000
bin_in=0110010001 bcd_out=0000010000000001
bin_in=0110010010 bcd_out=0000010000000010
bin_in=0110010011 bcd_out=0000010000000011
bin_in=0110010100 bcd_out=0000010000000100
bin_in=0110010101 bcd_out=0000010000000101
bin_in=0110010110 bcd_out=0000010000000110
bin_in=0110010111 bcd_out=0000010000000111
bin_in=0110011000 bcd_out=0000010000001000
bin_in=0110011001 bcd_out=0000010000001001
bin_in=0110011010 bcd_out=0000010000010000
bin_in=0110011011 bcd_out=0000010000010001
bin_in=0110011100 bcd_out=0000010000010010
bin_in=0110011101 bcd_out=0000010000010011
bin_in=0110011110 bcd_out=0000010000010100
bin_in=0110011111 bcd_out=0000010000010101
bin_in=0110100000 bcd_out=0000010000010110
bin_in=0110100001 bcd_out=0000010000010111
bin_in=0110100010 bcd_out=0000010000011000
bin_in=0110100011 bcd_out=0000010000011001
bin_in=0110100100 bcd_out=0000010000100000
bin_in=0110100101 bcd_out=0000010000100001
bin_in=0110100110 bcd_out=0000010000100010
bin_in=0110100111 bcd_out=0000010000100011
bin_in=0110101000 bcd_out=0000010000100100
bin_in=0110101001 bcd_out=0000010000100101
bin_in=0110101010 bcd_out=0000010000100110
bin_in=0110101011 bcd_out=0000010000100111
bin_in=0110101100 bcd_out=0000010000101000
bin_in=0110101101 bcd_out=0000010000101001
bin_in=0110101110 bcd_out=0000010000110000
bin_in=0110101111 bcd_out=0000010000110001
bin_in=0110110000 bcd_out=0000010000110010
bin_in=0110110001 bcd_out=0000010000110011
bin_in=0110110010 bcd_out=0000010000110100
bin_in=0110110011 bcd_out=0000010000110101
bin_in=0110110100 bcd_out=0000010000110110
bin_in=0110110101 bcd_out=0000010000110111
bin_in=0110110110 bcd_out=0000010000111000
bin_in=0110110111 bcd_out=0000010000111001
bin_in=0110111000 bcd_out=0000010001000000
bin_in=0110111001 bcd_out=0000010001000001
bin_in=0110111010 bcd_out=0000010001000010
bin_in=0110111011 bcd_out=0000010001000011
bin_in=0110111100 bcd_out=0000010001000100
bin_in=0110111101 bcd_out=0000010001000101
bin_in=0110111110 bcd_out=0000010001000110
bin_in=0110111111 bcd_out=0000010001000111
bin_in=0111000000 bcd_out=0000010001001000
bin_in=0111000001 bcd_out=0000010001001001
bin_in=0111000010 bcd_out=0000010001010000
bin_in=0111000011 bcd_out=0000010001010001
bin_in=0111000100 bcd_out=0000010001010010
bin_in=0111000101 bcd_out=0000010001010011
bin_in=0111000110 bcd_out=0000010001010100
bin_in=0111000111 bcd_out=0000010001010101
bin_in=0111001000 bcd_out=0000010001010110
bin_in=0111001001 bcd_out=0000010001010111
bin_in=0111001010 bcd_out=0000010001011000
bin_in=0111001011 bcd_out=0000010001011001
bin_in=0111001100 bcd_out=0000010001100000
bin_in=0111001101 bcd_out=0000010001100001
bin_in=0111001110 bcd_out=0000010001100010
bin_in=0111001111 bcd_out=0000010001100011
bin_in=0111010000 bcd_out=0000010001100100
bin_in=0111010001 bcd_out=0000010001100101
bin_in=0111010010 bcd_out=0000010001100110
bin_in=0111010011 bcd_out=0000010001100111
bin_in=0111010100 bcd_out=0000010001101000
bin_in=0111010101 bcd_out=0000010001101001
bin_in=0111010110 bcd_out=0000010001110000
bin_in=0111010111 bcd_out=0000010001110001
bin_in=0111011000 bcd_out=0000010001110010
bin_in=0111011001 bcd_out=0000010001110011
bin_in=0111011010 bcd_out=0000010001110100
bin_in=0111011011 bcd_out=0000010001110101
bin_in=0111011100 bcd_out=0000010001110110
bin_in=0111011101 bcd_out=0000010001110111
bin_in=0111011110 bcd_out=0000010001111000
bin_in=0111011111 bcd_out=0000010001111001
bin_in=0111100000 bcd_out=0000010010000000
bin_in=0111100001 bcd_out=0000010010000001
bin_in=0111100010 bcd_out=0000010010000010
bin_in=0111100011 bcd_out=0000010010000011
bin_in=0111100100 bcd_out=0000010010000100
bin_in=0111100101 bcd_out=0000010010000101
bin_in=0111100110 bcd_out=0000010010000110
bin_in=0111100111 bcd_out=0000010010000111
bin_in=0111101000 bcd_out=0000010010001000
bin_in=0111101001 bcd_out=0000010010001001
bin_in=0111101010 bcd_out=0000010010010000
bin_in=0111101011 bcd_out=0000010010010001
bin_in=0111101100 bcd_out=0000010010010010
bin_in=0111101101 bcd_out=0000010010010011
bin_in=0111101110 bcd_out=0000010010010100
bin_in=0111101111 bcd_out=0000010010010101
bin_in=0111110000 bcd_out=0000010010010110
bin_in=0111110001 bcd_out=0000010010010111
bin_in=0111110010 bcd_out=0000010010011000
bin_in=0111110011 bcd_out=0000010010011001
bin_in=0111110100 bcd_out=0000010100000000
bin_in=0111110101 bcd_out=0000010100000001
bin_in=0111110110 bcd_out=0000010100000010
bin_in=0111110111 bcd_out=0000010100000011
bin_in=0111111000 bcd_out=0000010100000100
bin_in=0111111001 bcd_out=0000010100000101
bin_in=0111111010 bcd_out=0000010100000110
bin_in=0111111011 bcd_out=0000010100000111
bin_in=0111111100 bcd_out=0000010100001000
bin_in=0111111101 bcd_out=0000010100001001
bin_in=0111111110 bcd_out=0000010100010000
bin_in=0111111111 bcd_out=0000010100010001
bin_in=1000000000 bcd_out=0000010100010010
bin_in=1000000001 bcd_out=0000010100010011
bin_in=1000000010 bcd_out=0000010100010100
bin_in=1000000011 bcd_out=0000010100010101
bin_in=1000000100 bcd_out=0000010100010110
bin_in=1000000101 bcd_out=0000010100010111
bin_in=1000000110 bcd_out=0000010100011000
bin_in=1000000111 bcd_out=0000010100011001
bin_in=1000001000 bcd_out=0000010100100000
bin_in=1000001001 bcd_out=0000010100100001
bin_in=1000001010 bcd_out=0000010100100010
bin_in=1000001011 bcd_out=0000010100100011
bin_in=1000001100 bcd_out=0000010100100100
bin_in=1000001101 bcd_out=0000010100100101
bin_in=1000001110 bcd_out=0000010100100110
bin_in=1000001111 bcd_out=0000010100100111
bin_in=1000010000 bcd_out=0000010100101000
bin_in=1000010001 bcd_out=0000010100101001
bin_in=1000010010 bcd_out=0000010100110000
bin_in=1000010011 bcd_out=0000010100110001
bin_in=1000010100 bcd_out=0000010100110010
bin_in=1000010101 bcd_out=0000010100110011
bin_in=1000010110 bcd_out=0000010100110100
bin_in=1000010111 bcd_out=0000010100110101
bin_in=1000011000 bcd_out=0000010100110110
bin_in=1000011001 bcd_out=0000010100110111
bin_in=1000011010 bcd_out=0000010100111000
bin_in=1000011011 bcd_out=0000010100111001
bin_in=1000011100 bcd_out=0000010101000000
bin_in=1000011101 bcd_out=0000010101000001
bin_in=1000011110 bcd_out=0000010101000010
bin_in=1000011111 bcd_out=0000010101000011
bin_in=1000100000 bcd_out=0000010101000100
bin_in=1000100001 bcd_out=0000010101000101
bin_in=1000100010 bcd_out=0000010101000110
bin_in=1000100011 bcd_out=0000010101000111
bin_in=1000100100 bcd_out=0000010101001000
bin_in=1000100101 bcd_out=0000010101001001
bin_in=1000100110 bcd_out=0000010101010000
bin_in=1000100111 bcd_out=0000010101010001
bin_in=1000101000 bcd_out=0000010101010010
bin_in=1000101001 bcd_out=0000010101010011
bin_in=1000101010 bcd_out=0000010101010100
bin_in=1000101011 bcd_out=0000010101010101
bin_in=1000101100 bcd_out=0000010101010110
bin_in=1000101101 bcd_out=0000010101010111
bin_in=1000101110 bcd_out=0000010101011000
bin_in=1000101111 bcd_out=0000010101011001
bin_in=1000110000 bcd_out=0000010101100000
bin_in=1000110001 bcd_out=0000010101100001
bin_in=1000110010 bcd_out=0000010101100010
bin_in=1000110011 bcd_out=0000010101100011
bin_in=1000110100 bcd_out=0000010101100100
bin_in=1000110101 bcd_out=0000010101100101
bin_in=1000110110 bcd_out=0000010101100110
bin_in=1000110111 bcd_out=0000010101100111
bin_in=1000111000 bcd_out=0000010101101000
bin_in=1000111001 bcd_out=0000010101101001
bin_in=1000111010 bcd_out=0000010101110000
bin_in=1000111011 bcd_out=0000010101110001
bin_in=1000111100 bcd_out=0000010101110010
bin_in=1000111101 bcd_out=0000010101110011
bin_in=1000111110 bcd_out=0000010101110100
bin_in=1000111111 bcd_out=0000010101110101
bin_in=1001000000 bcd_out=0000010101110110
bin_in=1001000001 bcd_out=0000010101110111
bin_in=1001000010 bcd_out=0000010101111000
bin_in=1001000011 bcd_out=0000010101111001
bin_in=1001000100 bcd_out=0000010110000000
bin_in=1001000101 bcd_out=0000010110000001
bin_in=1001000110 bcd_out=0000010110000010
bin_in=1001000111 bcd_out=0000010110000011
bin_in=1001001000 bcd_out=0000010110000100
bin_in=1001001001 bcd_out=0000010110000101
bin_in=1001001010 bcd_out=0000010110000110
bin_in=1001001011 bcd_out=0000010110000111
bin_in=1001001100 bcd_out=0000010110001000
bin_in=1001001101 bcd_out=0000010110001001
bin_in=1001001110 bcd_out=0000010110010000
bin_in=1001001111 bcd_out=0000010110010001
bin_in=1001010000 bcd_out=0000010110010010
bin_in=1001010001 bcd_out=0000010110010011
bin_in=1001010010 bcd_out=0000010110010100
bin_in=1001010011 bcd_out=0000010110010101
bin_in=1001010100 bcd_out=0000010110010110
bin_in=1001010101 bcd_out=0000010110010111
bin_in=1001010110 bcd_out=0000010110011000
bin_in=1001010111 bcd_out=0000010110011001
bin_in=1001011000 bcd_out=0000011000000000
bin_in=1001011001 bcd_out=0000011000000001
bin_in=1001011010 bcd_out=0000011000000010
bin_in=1001011011 bcd_out=0000011000000011
bin_in=1001011100 bcd_out=0000011000000100
bin_in=1001011101 bcd_out=0000011000000101
bin_in=1001011110 bcd_out=0000011000000110
bin_in=1001011111 bcd_out=0000011000000111
bin_in=1001100000 bcd_out=0000011000001000
bin_in=1001100001 bcd_out=0000011000001001
bin_in=1001100010 bcd_out=0000011000010000
bin_in=1001100011 bcd_out=0000011000010001
bin_in=1001100100 bcd_out=0000011000010010
bin_in=1001100101 bcd_out=0000011000010011
bin_in=1001100110 bcd_out=0000011000010100
bin_in=1001100111 bcd_out=0000011000010101
bin_in=1001101000 bcd_out=0000011000010110
bin_in=1001101001 bcd_out=0000011000010111
bin_in=1001101010 bcd_out=0000011000011000
bin_in=1001101011 bcd_out=0000011000011001
bin_in=1001101100 bcd_out=0000011000100000
bin_in=1001101101 bcd_out=0000011000100001
bin_in=1001101110 bcd_out=0000011000100010
bin_in=1001101111 bcd_out=0000011000100011
bin_in=1001110000 bcd_out=0000011000100100
bin_in=1001110001 bcd_out=0000011000100101
bin_in=1001110010 bcd_out=0000011000100110
bin_in=1001110011 bcd_out=0000011000100111
bin_in=1001110100 bcd_out=0000011000101000
bin_in=1001110101 bcd_out=0000011000101001
bin_in=1001110110 bcd_out=0000011000110000
bin_in=1001110111 bcd_out=0000011000110001
bin_in=1001111000 bcd_out=0000011000110010
bin_in=1001111001 bcd_out=0000011000110011
bin_in=1001111010 bcd_out=0000011000110100
bin_in=1001111011 bcd_out=0000011000110101
bin_in=1001111100 bcd_out=0000011000110110
bin_in=1001111101 bcd_out=0000011000110111
bin_in=1001111110 bcd_out=0000011000111000
bin_in=1001111111 bcd_out=0000011000111001
bin_in=1010000000 bcd_out=0000011001000000
bin_in=1010000001 bcd_out=0000011001000001
bin_in=1010000010 bcd_out=0000011001000010
bin_in=1010000011 bcd_out=0000011001000011
bin_in=1010000100 bcd_out=0000011001000100
bin_in=1010000101 bcd_out=0000011001000101
bin_in=1010000110 bcd_out=0000011001000110
bin_in=1010000111 bcd_out=0000011001000111
bin_in=1010001000 bcd_out=0000011001001000
bin_in=1010001001 bcd_out=0000011001001001
bin_in=1010001010 bcd_out=0000011001010000
bin_in=1010001011 bcd_out=0000011001010001
bin_in=1010001100 bcd_out=0000011001010010
bin_in=1010001101 bcd_out=0000011001010011
bin_in=1010001110 bcd_out=0000011001010100
bin_in=1010001111 bcd_out=0000011001010101
bin_in=1010010000 bcd_out=0000011001010110
bin_in=1010010001 bcd_out=0000011001010111
bin_in=1010010010 bcd_out=0000011001011000
bin_in=1010010011 bcd_out=0000011001011001
bin_in=1010010100 bcd_out=0000011001100000
bin_in=1010010101 bcd_out=0000011001100001
bin_in=1010010110 bcd_out=0000011001100010
bin_in=1010010111 bcd_out=0000011001100011
bin_in=1010011000 bcd_out=0000011001100100
bin_in=1010011001 bcd_out=0000011001100101
bin_in=1010011010 bcd_out=0000011001100110
bin_in=1010011011 bcd_out=0000011001100111
bin_in=1010011100 bcd_out=0000011001101000
bin_in=1010011101 bcd_out=0000011001101001
bin_in=1010011110 bcd_out=0000011001110000
bin_in=1010011111 bcd_out=0000011001110001
bin_in=1010100000 bcd_out=0000011001110010
bin_in=1010100001 bcd_out=0000011001110011
bin_in=1010100010 bcd_out=0000011001110100
bin_in=1010100011 bcd_out=0000011001110101
bin_in=1010100100 bcd_out=0000011001110110
bin_in=1010100101 bcd_out=0000011001110111
bin_in=1010100110 bcd_out=0000011001111000
bin_in=1010100111 bcd_out=0000011001111001
bin_in=1010101000 bcd_out=0000011010000000
bin_in=1010101001 bcd_out=0000011010000001
bin_in=1010101010 bcd_out=0000011010000010
bin_in=1010101011 bcd_out=0000011010000011
bin_in=1010101100 bcd_out=0000011010000100
bin_in=1010101101 bcd_out=0000011010000101
bin_in=1010101110 bcd_out=0000011010000110
bin_in=1010101111 bcd_out=0000011010000111
bin_in=1010110000 bcd_out=0000011010001000
bin_in=1010110001 bcd_out=0000011010001001
bin_in=1010110010 bcd_out=0000011010010000
bin_in=1010110011 bcd_out=0000011010010001
bin_in=1010110100 bcd_out=0000011010010010
bin_in=1010110101 bcd_out=0000011010010011
bin_in=1010110110 bcd_out=0000011010010100
bin_in=1010110111 bcd_out=0000011010010101
bin_in=1010111000 bcd_out=0000011010010110
bin_in=1010111001 bcd_out=0000011010010111
bin_in=1010111010 bcd_out=0000011010011000
bin_in=1010111011 bcd_out=0000011010011001
bin_in=1010111100 bcd_out=0000011100000000
bin_in=1010111101 bcd_out=0000011100000001
bin_in=1010111110 bcd_out=0000011100000010
bin_in=1010111111 bcd_out=0000011100000011
bin_in=1011000000 bcd_out=0000011100000100
bin_in=1011000001 bcd_out=0000011100000101
bin_in=1011000010 bcd_out=0000011100000110
bin_in=1011000011 bcd_out=0000011100000111
bin_in=1011000100 bcd_out=0000011100001000
bin_in=1011000101 bcd_out=0000011100001001
bin_in=1011000110 bcd_out=0000011100010000
bin_in=1011000111 bcd_out=0000011100010001
bin_in=1011001000 bcd_out=0000011100010010
bin_in=1011001001 bcd_out=0000011100010011
bin_in=1011001010 bcd_out=0000011100010100
bin_in=1011001011 bcd_out=0000011100010101
bin_in=1011001100 bcd_out=0000011100010110
bin_in=1011001101 bcd_out=0000011100010111
bin_in=1011001110 bcd_out=0000011100011000
bin_in=1011001111 bcd_out=0000011100011001
bin_in=1011010000 bcd_out=0000011100100000
bin_in=1011010001 bcd_out=0000011100100001
bin_in=1011010010 bcd_out=0000011100100010
bin_in=1011010011 bcd_out=0000011100100011
bin_in=1011010100 bcd_out=0000011100100100
bin_in=1011010101 bcd_out=0000011100100101
bin_in=1011010110 bcd_out=0000011100100110
bin_in=1011010111 bcd_out=0000011100100111
bin_in=1011011000 bcd_out=0000011100101000
bin_in=1011011001 bcd_out=0000011100101001
bin_in=1011011010 bcd_out=0000011100110000
bin_in=1011011011 bcd_out=0000011100110001
bin_in=1011011100 bcd_out=0000011100110010
bin_in=1011011101 bcd_out=0000011100110011
bin_in=1011011110 bcd_out=0000011100110100
bin_in=1011011111 bcd_out=0000011100110101
bin_in=1011100000 bcd_out=0000011100110110
bin_in=1011100001 bcd_out=0000011100110111
bin_in=1011100010 bcd_out=0000011100111000
bin_in=1011100011 bcd_out=0000011100111001
bin_in=1011100100 bcd_out=0000011101000000
bin_in=1011100101 bcd_out=0000011101000001
bin_in=1011100110 bcd_out=0000011101000010
bin_in=1011100111 bcd_out=0000011101000011
bin_in=1011101000 bcd_out=0000011101000100
bin_in=1011101001 bcd_out=0000011101000101
bin_in=1011101010 bcd_out=0000011101000110
bin_in=1011101011 bcd_out=0000011101000111
bin_in=1011101100 bcd_out=0000011101001000
bin_in=1011101101 bcd_out=0000011101001001
bin_in=1011101110 bcd_out=0000011101010000
bin_in=1011101111 bcd_out=0000011101010001
bin_in=1011110000 bcd_out=0000011101010010
bin_in=1011110001 bcd_out=0000011101010011
bin_in=1011110010 bcd_out=0000011101010100
bin_in=1011110011 bcd_out=0000011101010101
bin_in=1011110100 bcd_out=0000011101010110
bin_in=1011110101 bcd_out=0000011101010111
bin_in=1011110110 bcd_out=0000011101011000
bin_in=1011110111 bcd_out=0000011101011001
bin_in=1011111000 bcd_out=0000011101100000
bin_in=1011111001 bcd_out=0000011101100001
bin_in=1011111010 bcd_out=0000011101100010
bin_in=1011111011 bcd_out=0000011101100011
bin_in=1011111100 bcd_out=0000011101100100
bin_in=1011111101 bcd_out=0000011101100101
bin_in=1011111110 bcd_out=0000011101100110
bin_in=1011111111 bcd_out=0000011101100111
bin_in=1100000000 bcd_out=0000011101101000
bin_in=1100000001 bcd_out=0000011101101001
bin_in=1100000010 bcd_out=0000011101110000
bin_in=1100000011 bcd_out=0000011101110001
bin_in=1100000100 bcd_out=0000011101110010
bin_in=1100000101 bcd_out=0000011101110011
bin_in=1100000110 bcd_out=0000011101110100
bin_in=1100000111 bcd_out=0000011101110101
bin_in=1100001000 bcd_out=0000011101110110
bin_in=1100001001 bcd_out=0000011101110111
bin_in=1100001010 bcd_out=0000011101111000
bin_in=1100001011 bcd_out=0000011101111001
bin_in=1100001100 bcd_out=0000011110000000
bin_in=1100001101 bcd_out=0000011110000001
bin_in=1100001110 bcd_out=0000011110000010
bin_in=1100001111 bcd_out=0000011110000011
bin_in=1100010000 bcd_out=0000011110000100
bin_in=1100010001 bcd_out=0000011110000101
bin_in=1100010010 bcd_out=0000011110000110
bin_in=1100010011 bcd_out=0000011110000111
bin_in=1100010100 bcd_out=0000011110001000
bin_in=1100010101 bcd_out=0000011110001001
bin_in=1100010110 bcd_out=0000011110010000
bin_in=1100010111 bcd_out=0000011110010001
bin_in=1100011000 bcd_out=0000011110010010
bin_in=1100011001 bcd_out=0000011110010011
bin_in=1100011010 bcd_out=0000011110010100
bin_in=1100011011 bcd_out=0000011110010101
bin_in=1100011100 bcd_out=0000011110010110
bin_in=1100011101 bcd_out=0000011110010111
bin_in=1100011110 bcd_out=0000011110011000
bin_in=1100011111 bcd_out=0000011110011001
bin_in=1100100000 bcd_out=0000100000000000
bin_in=1100100001 bcd_out=0000100000000001
bin_in=1100100010 bcd_out=0000100000000010
bin_in=1100100011 bcd_out=0000100000000011
bin_in=1100100100 bcd_out=0000100000000100
bin_in=1100100101 bcd_out=0000100000000101
bin_in=1100100110 bcd_out=0000100000000110
bin_in=1100100111 bcd_out=0000100000000111
bin_in=1100101000 bcd_out=0000100000001000
bin_in=1100101001 bcd_out=0000100000001001
bin_in=1100101010 bcd_out=0000100000010000
bin_in=1100101011 bcd_out=0000100000010001
bin_in=1100101100 bcd_out=0000100000010010
bin_in=1100101101 bcd_out=0000100000010011
bin_in=1100101110 bcd_out=0000100000010100
bin_in=1100101111 bcd_out=0000100000010101
bin_in=1100110000 bcd_out=0000100000010110
bin_in=1100110001 bcd_out=0000100000010111
bin_in=1100110010 bcd_out=0000100000011000
bin_in=1100110011 bcd_out=0000100000011001
bin_in=1100110100 bcd_out=0000100000100000
bin_in=1100110101 bcd_out=0000100000100001
bin_in=1100110110 bcd_out=0000100000100010
bin_in=1100110111 bcd_out=0000100000100011
bin_in=1100111000 bcd_out=0000100000100100
bin_in=1100111001 bcd_out=0000100000100101
bin_in=1100111010 bcd_out=0000100000100110
bin_in=1100111011 bcd_out=0000100000100111
bin_in=1100111100 bcd_out=0000100000101000
bin_in=1100111101 bcd_out=0000100000101001
bin_in=1100111110 bcd_out=0000100000110000
bin_in=1100111111 bcd_out=0000100000110001
bin_in=1101000000 bcd_out=0000100000110010
bin_in=1101000001 bcd_out=0000100000110011
bin_in=1101000010 bcd_out=0000100000110100
bin_in=1101000011 bcd_out=0000100000110101
bin_in=1101000100 bcd_out=0000100000110110
bin_in=1101000101 bcd_out=0000100000110111
bin_in=1101000110 bcd_out=0000100000111000
bin_in=1101000111 bcd_out=0000100000111001
bin_in=1101001000 bcd_out=0000100001000000
bin_in=1101001001 bcd_out=0000100001000001
bin_in=1101001010 bcd_out=0000100001000010
bin_in=1101001011 bcd_out=0000100001000011
bin_in=1101001100 bcd_out=0000100001000100
bin_in=1101001101 bcd_out=0000100001000101
bin_in=1101001110 bcd_out=0000100001000110
bin_in=1101001111 bcd_out=0000100001000111
bin_in=1101010000 bcd_out=0000100001001000
bin_in=1101010001 bcd_out=0000100001001001
bin_in=1101010010 bcd_out=0000100001010000
bin_in=1101010011 bcd_out=0000100001010001
bin_in=1101010100 bcd_out=0000100001010010
bin_in=1101010101 bcd_out=0000100001010011
bin_in=1101010110 bcd_out=0000100001010100
bin_in=1101010111 bcd_out=0000100001010101
bin_in=1101011000 bcd_out=0000100001010110
bin_in=1101011001 bcd_out=0000100001010111
bin_in=1101011010 bcd_out=0000100001011000
bin_in=1101011011 bcd_out=0000100001011001
bin_in=1101011100 bcd_out=0000100001100000
bin_in=1101011101 bcd_out=0000100001100001
bin_in=1101011110 bcd_out=0000100001100010
bin_in=1101011111 bcd_out=0000100001100011
bin_in=1101100000 bcd_out=0000100001100100
bin_in=1101100001 bcd_out=0000100001100101
bin_in=1101100010 bcd_out=0000100001100110
bin_in=1101100011 bcd_out=0000100001100111
bin_in=1101100100 bcd_out=0000100001101000
bin_in=1101100101 bcd_out=0000100001101001
bin_in=1101100110 bcd_out=0000100001110000
bin_in=1101100111 bcd_out=0000100001110001
bin_in=1101101000 bcd_out=0000100001110010
bin_in=1101101001 bcd_out=0000100001110011
bin_in=1101101010 bcd_out=0000100001110100
bin_in=1101101011 bcd_out=0000100001110101
bin_in=1101101100 bcd_out=0000100001110110
bin_in=1101101101 bcd_out=0000100001110111
bin_in=1101101110 bcd_out=0000100001111000
bin_in=1101101111 bcd_out=0000100001111001
bin_in=1101110000 bcd_out=0000100010000000
bin_in=1101110001 bcd_out=0000100010000001
bin_in=1101110010 bcd_out=0000100010000010
bin_in=1101110011 bcd_out=0000100010000011
bin_in=1101110100 bcd_out=0000100010000100
bin_in=1101110101 bcd_out=0000100010000101
bin_in=1101110110 bcd_out=0000100010000110
bin_in=1101110111 bcd_out=0000100010000111
bin_in=1101111000 bcd_out=0000100010001000
bin_in=1101111001 bcd_out=0000100010001001
bin_in=1101111010 bcd_out=0000100010010000
bin_in=1101111011 bcd_out=0000100010010001
bin_in=1101111100 bcd_out=0000100010010010
bin_in=1101111101 bcd_out=0000100010010011
bin_in=1101111110 bcd_out=0000100010010100
bin_in=1101111111 bcd_out=0000100010010101
bin_in=1110000000 bcd_out=0000100010010110
bin_in=1110000001 bcd_out=0000100010010111
bin_in=1110000010 bcd_out=0000100010011000
bin_in=1110000011 bcd_out=0000100010011001
bin_in=1110000100 bcd_out=0000100100000000
bin_in=1110000101 bcd_out=0000100100000001
bin_in=1110000110 bcd_out=0000100100000010
bin_in=1110000111 bcd_out=0000100100000011
bin_in=1110001000 bcd_out=0000100100000100
bin_in=1110001001 bcd_out=0000100100000101
bin_in=1110001010 bcd_out=0000100100000110
bin_in=1110001011 bcd_out=0000100100000111
bin_in=1110001100 bcd_out=0000100100001000
bin_in=1110001101 bcd_out=0000100100001001
bin_in=1110001110 bcd_out=0000100100010000
bin_in=1110001111 bcd_out=0000100100010001
bin_in=1110010000 bcd_out=0000100100010010
bin_in=1110010001 bcd_out=0000100100010011
bin_in=1110010010 bcd_out=0000100100010100
bin_in=1110010011 bcd_out=0000100100010101
bin_in=1110010100 bcd_out=0000100100010110
bin_in=1110010101 bcd_out=0000100100010111
bin_in=1110010110 bcd_out=0000100100011000
bin_in=1110010111 bcd_out=0000100100011001
bin_in=1110011000 bcd_out=0000100100100000
bin_in=1110011001 bcd_out=0000100100100001
bin_in=1110011010 bcd_out=0000100100100010
bin_in=1110011011 bcd_out=0000100100100011
bin_in=1110011100 bcd_out=0000100100100100
bin_in=1110011101 bcd_out=0000100100100101
bin_in=1110011110 bcd_out=0000100100100110
bin_in=1110011111 bcd_out=0000100100100111
bin_in=1110100000 bcd_out=0000100100101000
bin_in=1110100001 bcd_out=0000100100101001
bin_in=1110100010 bcd_out=0000100100110000
bin_in=1110100011 bcd_out=0000100100110001
bin_in=1110100100 bcd_out=0000100100110010
bin_in=1110100101 bcd_out=0000100100110011
bin_in=1110100110 bcd_out=0000100100110100
bin_in=1110100111 bcd_out=0000100100110101
bin_in=1110101000 bcd_out=0000100100110110
bin_in=1110101001 bcd_out=0000100100110111
bin_in=1110101010 bcd_out=0000100100111000
bin_in=1110101011 bcd_out=0000100100111001
bin_in=1110101100 bcd_out=0000100101000000
bin_in=1110101101 bcd_out=0000100101000001
bin_in=1110101110 bcd_out=0000100101000010
bin_in=1110101111 bcd_out=0000100101000011
bin_in=1110110000 bcd_out=0000100101000100
bin_in=1110110001 bcd_out=0000100101000101
bin_in=1110110010 bcd_out=0000100101000110
bin_in=1110110011 bcd_out=0000100101000111
bin_in=1110110100 bcd_out=0000100101001000
bin_in=1110110101 bcd_out=0000100101001001
bin_in=1110110110 bcd_out=0000100101010000
bin_in=1110110111 bcd_out=0000100101010001
bin_in=1110111000 bcd_out=0000100101010010
bin_in=1110111001 bcd_out=0000100101010011
bin_in=1110111010 bcd_out=0000100101010100
bin_in=1110111011 bcd_out=0000100101010101
bin_in=1110111100 bcd_out=0000100101010110
bin_in=1110111101 bcd_out=0000100101010111
bin_in=1110111110 bcd_out=0000100101011000
bin_in=1110111111 bcd_out=0000100101011001
bin_in=1111000000 bcd_out=0000100101100000
bin_in=1111000001 bcd_out=0000100101100001
bin_in=1111000010 bcd_out=0000100101100010
bin_in=1111000011 bcd_out=0000100101100011
bin_in=1111000100 bcd_out=0000100101100100
bin_in=1111000101 bcd_out=0000100101100101
bin_in=1111000110 bcd_out=0000100101100110
bin_in=1111000111 bcd_out=0000100101100111
bin_in=1111001000 bcd_out=0000100101101000
bin_in=1111001001 bcd_out=0000100101101001
bin_in=1111001010 bcd_out=0000100101110000
bin_in=1111001011 bcd_out=0000100101110001
bin_in=1111001100 bcd_out=0000100101110010
bin_in=1111001101 bcd_out=0000100101110011
bin_in=1111001110 bcd_out=0000100101110100
bin_in=1111001111 bcd_out=0000100101110101
bin_in=1111010000 bcd_out=0000100101110110
bin_in=1111010001 bcd_out=0000100101110111
bin_in=1111010010 bcd_out=0000100101111000
bin_in=1111010011 bcd_out=0000100101111001
bin_in=1111010100 bcd_out=0000100110000000
bin_in=1111010101 bcd_out=0000100110000001
bin_in=1111010110 bcd_out=0000100110000010
bin_in=1111010111 bcd_out=0000100110000011
bin_in=1111011000 bcd_out=0000100110000100
bin_in=1111011001 bcd_out=0000100110000101
bin_in=1111011010 bcd_out=0000100110000110
bin_in=1111011011 bcd_out=0000100110000111
bin_in=1111011100 bcd_out=0000100110001000
bin_in=1111011101 bcd_out=0000100110001001
bin_in=1111011110 bcd_out=0000100110010000
bin_in=1111011111 bcd_out=0000100110010001
bin_in=1111100000 bcd_out=0000100110010010
bin_in=1111100001 bcd_out=0000100110010011
bin_in=1111100010 bcd_out=0000100110010100
bin_in=1111100011 bcd_out=0000100110010101
bin_in=1111100100 bcd_out=0000100110010110
bin_in=1111100101 bcd_out=0000100110010111
bin_in=1111100110 bcd_out=0000100110011000
bin_in=1111100111 bcd_out=0000100110011001
bin_in=1111101000 bcd_out=0001000000000000
bin_in=1111101001 bcd_out=0001000000000001
bin_in=1111101010 bcd_out=0001000000000010
bin_in=1111101011 bcd_out=0001000000000011
bin_in=1111101100 bcd_out=0001000000000100
bin_in=1111101101 bcd_out=0001000000000101
bin_in=1111101110 bcd_out=0001000000000110
bin_in=1111101111 bcd_out=0001000000000111
bin_in=1111110000 bcd_out=0001000000001000
bin_in=1111110001 bcd_out=0001000000001001
bin_in=1111110010 bcd_out=0001000000010000
bin_in=1111110011 bcd_out=0001000000010001
bin_in=1111110100 bcd_out=0001000000010010
bin_in=1111110101 bcd_out=0001000000010011
bin_in=1111110110 bcd_out=0001000000010100
bin_in=1111110111 bcd_out=0001000000010101
bin_in=1111111000 bcd_out=0001000000010110
bin_in=1111111001 bcd_out=0001000000010111
bin_in=1111111010 bcd_out=0001000000011000
bin_in=1111111011 bcd_out=0001000000011001
bin_in=1111111100 bcd_out=0001000000100000
bin_in=1111111101 bcd_out=0001000000100001
bin_in=1111111110 bcd_out=0001000000100010
bin_in=1111111111 bcd_out=0001000000100011
binary_to_bcd_tb.v:20: $finish called at 10240 (1s)
* 
*/
